module spi_mvp(
    input clk100m,
    input rst,

    input sck,
    output miso,
    input mosi,
    input ss,

);

endmodule
