// Polyphase filter bank for upsampling from 44100.0kHz to 48000.0kHz
// Depth: 32

module rom_firbank_441_480(
    input clk,
    input [11:0] addr,
    output [23:0] data);
reg [23:0] data_ff;
assign data = data_ff;
always @(posedge clk) begin
    case(addr)
        0: data_ff <= 24'd44320;
        1: data_ff <= -24'd29396;
        2: data_ff <= 24'd22678;
        3: data_ff <= -24'd17801;
        4: data_ff <= 24'd13701;
        5: data_ff <= -24'd10175;
        6: data_ff <= 24'd7217;
        7: data_ff <= -24'd4849;
        8: data_ff <= 24'd3058;
        9: data_ff <= -24'd1790;
        10: data_ff <= 24'd959;
        11: data_ff <= -24'd460;
        12: data_ff <= 24'd191;
        13: data_ff <= -24'd63;
        14: data_ff <= 24'd13;
        15: data_ff <= -24'd1;
        16: data_ff <= 24'd96251;
        17: data_ff <= -24'd53535;
        18: data_ff <= 24'd37032;
        19: data_ff <= -24'd26973;
        20: data_ff <= 24'd19658;
        21: data_ff <= -24'd14003;
        22: data_ff <= 24'd9612;
        23: data_ff <= -24'd6289;
        24: data_ff <= 24'd3881;
        25: data_ff <= -24'd2231;
        26: data_ff <= 24'd1177;
        27: data_ff <= -24'd557;
        28: data_ff <= 24'd229;
        29: data_ff <= -24'd75;
        30: data_ff <= 24'd16;
        31: data_ff <= -24'd1;
        32: data_ff <= 24'd148834;
        33: data_ff <= -24'd77832;
        34: data_ff <= 24'd51456;
        35: data_ff <= -24'd36185;
        36: data_ff <= 24'd25639;
        37: data_ff <= -24'd17847;
        38: data_ff <= 24'd12018;
        39: data_ff <= -24'd7736;
        40: data_ff <= 24'd4708;
        41: data_ff <= -24'd2675;
        42: data_ff <= 24'd1397;
        43: data_ff <= -24'd656;
        44: data_ff <= 24'd267;
        45: data_ff <= -24'd87;
        46: data_ff <= 24'd18;
        47: data_ff <= -24'd1;
        48: data_ff <= 24'd202059;
        49: data_ff <= -24'd102279;
        50: data_ff <= 24'd65945;
        51: data_ff <= -24'd45433;
        52: data_ff <= 24'd31643;
        53: data_ff <= -24'd21707;
        54: data_ff <= 24'd14433;
        55: data_ff <= -24'd9190;
        56: data_ff <= 24'd5540;
        57: data_ff <= -24'd3121;
        58: data_ff <= 24'd1618;
        59: data_ff <= -24'd755;
        60: data_ff <= 24'd305;
        61: data_ff <= -24'd100;
        62: data_ff <= 24'd21;
        63: data_ff <= -24'd1;
        64: data_ff <= 24'd255920;
        65: data_ff <= -24'd126869;
        66: data_ff <= 24'd80494;
        67: data_ff <= -24'd54713;
        68: data_ff <= 24'd37667;
        69: data_ff <= -24'd25579;
        70: data_ff <= 24'd16858;
        71: data_ff <= -24'd10650;
        72: data_ff <= 24'd6375;
        73: data_ff <= -24'd3570;
        74: data_ff <= 24'd1841;
        75: data_ff <= -24'd854;
        76: data_ff <= 24'd344;
        77: data_ff <= -24'd112;
        78: data_ff <= 24'd23;
        79: data_ff <= -24'd2;
        80: data_ff <= 24'd310407;
        81: data_ff <= -24'd151593;
        82: data_ff <= 24'd95097;
        83: data_ff <= -24'd64022;
        84: data_ff <= 24'd43710;
        85: data_ff <= -24'd29464;
        86: data_ff <= 24'd19291;
        87: data_ff <= -24'd12116;
        88: data_ff <= 24'd7214;
        89: data_ff <= -24'd4021;
        90: data_ff <= 24'd2064;
        91: data_ff <= -24'd955;
        92: data_ff <= 24'd384;
        93: data_ff <= -24'd125;
        94: data_ff <= 24'd26;
        95: data_ff <= -24'd2;
        96: data_ff <= 24'd365512;
        97: data_ff <= -24'd176443;
        98: data_ff <= 24'd109749;
        99: data_ff <= -24'd73357;
        100: data_ff <= 24'd49768;
        101: data_ff <= -24'd33359;
        102: data_ff <= 24'd21731;
        103: data_ff <= -24'd13586;
        104: data_ff <= 24'd8057;
        105: data_ff <= -24'd4474;
        106: data_ff <= 24'd2290;
        107: data_ff <= -24'd1056;
        108: data_ff <= 24'd424;
        109: data_ff <= -24'd138;
        110: data_ff <= 24'd29;
        111: data_ff <= -24'd2;
        112: data_ff <= 24'd421227;
        113: data_ff <= -24'd201411;
        114: data_ff <= 24'd124446;
        115: data_ff <= -24'd82714;
        116: data_ff <= 24'd55839;
        117: data_ff <= -24'd37263;
        118: data_ff <= 24'd24178;
        119: data_ff <= -24'd15061;
        120: data_ff <= 24'd8902;
        121: data_ff <= -24'd4929;
        122: data_ff <= 24'd2516;
        123: data_ff <= -24'd1158;
        124: data_ff <= 24'd464;
        125: data_ff <= -24'd150;
        126: data_ff <= 24'd32;
        127: data_ff <= -24'd2;
        128: data_ff <= 24'd477542;
        129: data_ff <= -24'd226488;
        130: data_ff <= 24'd139181;
        131: data_ff <= -24'd92090;
        132: data_ff <= 24'd61921;
        133: data_ff <= -24'd41175;
        134: data_ff <= 24'd26630;
        135: data_ff <= -24'd16540;
        136: data_ff <= 24'd9750;
        137: data_ff <= -24'd5386;
        138: data_ff <= 24'd2743;
        139: data_ff <= -24'd1260;
        140: data_ff <= 24'd504;
        141: data_ff <= -24'd164;
        142: data_ff <= 24'd34;
        143: data_ff <= -24'd2;
        144: data_ff <= 24'd534449;
        145: data_ff <= -24'd251665;
        146: data_ff <= 24'd153948;
        147: data_ff <= -24'd101481;
        148: data_ff <= 24'd68013;
        149: data_ff <= -24'd45093;
        150: data_ff <= 24'd29086;
        151: data_ff <= -24'd18022;
        152: data_ff <= 24'd10601;
        153: data_ff <= -24'd5844;
        154: data_ff <= 24'd2972;
        155: data_ff <= -24'd1363;
        156: data_ff <= 24'd545;
        157: data_ff <= -24'd177;
        158: data_ff <= 24'd37;
        159: data_ff <= -24'd3;
        160: data_ff <= 24'd591938;
        161: data_ff <= -24'd276935;
        162: data_ff <= 24'd168744;
        163: data_ff <= -24'd110883;
        164: data_ff <= 24'd74110;
        165: data_ff <= -24'd49015;
        166: data_ff <= 24'd31545;
        167: data_ff <= -24'd19507;
        168: data_ff <= 24'd11454;
        169: data_ff <= -24'd6304;
        170: data_ff <= 24'd3201;
        171: data_ff <= -24'd1467;
        172: data_ff <= 24'd586;
        173: data_ff <= -24'd190;
        174: data_ff <= 24'd40;
        175: data_ff <= -24'd3;
        176: data_ff <= 24'd650000;
        177: data_ff <= -24'd302288;
        178: data_ff <= 24'd183561;
        179: data_ff <= -24'd120294;
        180: data_ff <= 24'd80212;
        181: data_ff <= -24'd52940;
        182: data_ff <= 24'd34008;
        183: data_ff <= -24'd20993;
        184: data_ff <= 24'd12308;
        185: data_ff <= -24'd6765;
        186: data_ff <= 24'd3431;
        187: data_ff <= -24'd1571;
        188: data_ff <= 24'd627;
        189: data_ff <= -24'd203;
        190: data_ff <= 24'd43;
        191: data_ff <= -24'd3;
        192: data_ff <= 24'd708625;
        193: data_ff <= -24'd327715;
        194: data_ff <= 24'd198394;
        195: data_ff <= -24'd129708;
        196: data_ff <= 24'd86315;
        197: data_ff <= -24'd56866;
        198: data_ff <= 24'd36471;
        199: data_ff <= -24'd22482;
        200: data_ff <= 24'd13164;
        201: data_ff <= -24'd7228;
        202: data_ff <= 24'd3662;
        203: data_ff <= -24'd1676;
        204: data_ff <= 24'd668;
        205: data_ff <= -24'd217;
        206: data_ff <= 24'd46;
        207: data_ff <= -24'd3;
        208: data_ff <= 24'd767803;
        209: data_ff <= -24'd353208;
        210: data_ff <= 24'd213239;
        211: data_ff <= -24'd139123;
        212: data_ff <= 24'd92418;
        213: data_ff <= -24'd60793;
        214: data_ff <= 24'd38936;
        215: data_ff <= -24'd23971;
        216: data_ff <= 24'd14020;
        217: data_ff <= -24'd7691;
        218: data_ff <= 24'd3894;
        219: data_ff <= -24'd1781;
        220: data_ff <= 24'd710;
        221: data_ff <= -24'd231;
        222: data_ff <= 24'd49;
        223: data_ff <= -24'd3;
        224: data_ff <= 24'd827525;
        225: data_ff <= -24'd378757;
        226: data_ff <= 24'd228088;
        227: data_ff <= -24'd148535;
        228: data_ff <= 24'd98517;
        229: data_ff <= -24'd64717;
        230: data_ff <= 24'd41399;
        231: data_ff <= -24'd25461;
        232: data_ff <= 24'd14878;
        233: data_ff <= -24'd8154;
        234: data_ff <= 24'd4126;
        235: data_ff <= -24'd1886;
        236: data_ff <= 24'd752;
        237: data_ff <= -24'd245;
        238: data_ff <= 24'd53;
        239: data_ff <= -24'd4;
        240: data_ff <= 24'd887780;
        241: data_ff <= -24'd404354;
        242: data_ff <= 24'd242937;
        243: data_ff <= -24'd157940;
        244: data_ff <= 24'd104611;
        245: data_ff <= -24'd68639;
        246: data_ff <= 24'd43862;
        247: data_ff <= -24'd26950;
        248: data_ff <= 24'd15735;
        249: data_ff <= -24'd8619;
        250: data_ff <= 24'd4359;
        251: data_ff <= -24'd1992;
        252: data_ff <= 24'd794;
        253: data_ff <= -24'd258;
        254: data_ff <= 24'd56;
        255: data_ff <= -24'd4;
        256: data_ff <= 24'd948557;
        257: data_ff <= -24'd429989;
        258: data_ff <= 24'd257780;
        259: data_ff <= -24'd167335;
        260: data_ff <= 24'd110697;
        261: data_ff <= -24'd72555;
        262: data_ff <= 24'd46322;
        263: data_ff <= -24'd28439;
        264: data_ff <= 24'd16593;
        265: data_ff <= -24'd9083;
        266: data_ff <= 24'd4592;
        267: data_ff <= -24'd2098;
        268: data_ff <= 24'd837;
        269: data_ff <= -24'd272;
        270: data_ff <= 24'd59;
        271: data_ff <= -24'd4;
        272: data_ff <= 24'd1009847;
        273: data_ff <= -24'd455653;
        274: data_ff <= 24'd272610;
        275: data_ff <= -24'd176715;
        276: data_ff <= 24'd116773;
        277: data_ff <= -24'd76466;
        278: data_ff <= 24'd48779;
        279: data_ff <= -24'd29926;
        280: data_ff <= 24'd17450;
        281: data_ff <= -24'd9548;
        282: data_ff <= 24'd4825;
        283: data_ff <= -24'd2204;
        284: data_ff <= 24'd879;
        285: data_ff <= -24'd287;
        286: data_ff <= 24'd62;
        287: data_ff <= -24'd4;
        288: data_ff <= 24'd1071638;
        289: data_ff <= -24'd481336;
        290: data_ff <= 24'd287423;
        291: data_ff <= -24'd186078;
        292: data_ff <= 24'd122836;
        293: data_ff <= -24'd80368;
        294: data_ff <= 24'd51231;
        295: data_ff <= -24'd31411;
        296: data_ff <= 24'd18307;
        297: data_ff <= -24'd10013;
        298: data_ff <= 24'd5059;
        299: data_ff <= -24'd2311;
        300: data_ff <= 24'd922;
        301: data_ff <= -24'd301;
        302: data_ff <= 24'd66;
        303: data_ff <= -24'd5;
        304: data_ff <= 24'd1133920;
        305: data_ff <= -24'd507030;
        306: data_ff <= 24'd302211;
        307: data_ff <= -24'd195419;
        308: data_ff <= 24'd128883;
        309: data_ff <= -24'd84260;
        310: data_ff <= 24'd53678;
        311: data_ff <= -24'd32894;
        312: data_ff <= 24'd19162;
        313: data_ff <= -24'd10477;
        314: data_ff <= 24'd5293;
        315: data_ff <= -24'd2417;
        316: data_ff <= 24'd965;
        317: data_ff <= -24'd315;
        318: data_ff <= 24'd69;
        319: data_ff <= -24'd5;
        320: data_ff <= 24'd1196681;
        321: data_ff <= -24'd532725;
        322: data_ff <= 24'd316971;
        323: data_ff <= -24'd204734;
        324: data_ff <= 24'd134913;
        325: data_ff <= -24'd88142;
        326: data_ff <= 24'd56118;
        327: data_ff <= -24'd34373;
        328: data_ff <= 24'd20017;
        329: data_ff <= -24'd10941;
        330: data_ff <= 24'd5526;
        331: data_ff <= -24'd2524;
        332: data_ff <= 24'd1008;
        333: data_ff <= -24'd329;
        334: data_ff <= 24'd72;
        335: data_ff <= -24'd5;
        336: data_ff <= 24'd1259911;
        337: data_ff <= -24'd558410;
        338: data_ff <= 24'd331695;
        339: data_ff <= -24'd214020;
        340: data_ff <= 24'd140923;
        341: data_ff <= -24'd92011;
        342: data_ff <= 24'd58552;
        343: data_ff <= -24'd35848;
        344: data_ff <= 24'd20869;
        345: data_ff <= -24'd11405;
        346: data_ff <= 24'd5760;
        347: data_ff <= -24'd2631;
        348: data_ff <= 24'd1051;
        349: data_ff <= -24'd344;
        350: data_ff <= 24'd76;
        351: data_ff <= -24'd5;
        352: data_ff <= 24'd1323597;
        353: data_ff <= -24'd584078;
        354: data_ff <= 24'd346377;
        355: data_ff <= -24'd223273;
        356: data_ff <= 24'd146909;
        357: data_ff <= -24'd95865;
        358: data_ff <= 24'd60976;
        359: data_ff <= -24'd37319;
        360: data_ff <= 24'd21719;
        361: data_ff <= -24'd11868;
        362: data_ff <= 24'd5993;
        363: data_ff <= -24'd2738;
        364: data_ff <= 24'd1094;
        365: data_ff <= -24'd358;
        366: data_ff <= 24'd79;
        367: data_ff <= -24'd6;
        368: data_ff <= 24'd1387729;
        369: data_ff <= -24'd609717;
        370: data_ff <= 24'd361013;
        371: data_ff <= -24'd232490;
        372: data_ff <= 24'd152871;
        373: data_ff <= -24'd99704;
        374: data_ff <= 24'd63392;
        375: data_ff <= -24'd38785;
        376: data_ff <= 24'd22567;
        377: data_ff <= -24'd12329;
        378: data_ff <= 24'd6226;
        379: data_ff <= -24'd2845;
        380: data_ff <= 24'd1138;
        381: data_ff <= -24'd373;
        382: data_ff <= 24'd83;
        383: data_ff <= -24'd6;
        384: data_ff <= 24'd1452294;
        385: data_ff <= -24'd635318;
        386: data_ff <= 24'd375595;
        387: data_ff <= -24'd241665;
        388: data_ff <= 24'd158805;
        389: data_ff <= -24'd103524;
        390: data_ff <= 24'd65796;
        391: data_ff <= -24'd40245;
        392: data_ff <= 24'd23412;
        393: data_ff <= -24'd12790;
        394: data_ff <= 24'd6459;
        395: data_ff <= -24'd2952;
        396: data_ff <= 24'd1181;
        397: data_ff <= -24'd388;
        398: data_ff <= 24'd86;
        399: data_ff <= -24'd6;
        400: data_ff <= 24'd1517281;
        401: data_ff <= -24'd660871;
        402: data_ff <= 24'd390119;
        403: data_ff <= -24'd250797;
        404: data_ff <= 24'd164709;
        405: data_ff <= -24'd107326;
        406: data_ff <= 24'd68190;
        407: data_ff <= -24'd41698;
        408: data_ff <= 24'd24254;
        409: data_ff <= -24'd13249;
        410: data_ff <= 24'd6691;
        411: data_ff <= -24'd3059;
        412: data_ff <= 24'd1224;
        413: data_ff <= -24'd402;
        414: data_ff <= 24'd90;
        415: data_ff <= -24'd7;
        416: data_ff <= 24'd1582678;
        417: data_ff <= -24'd686367;
        418: data_ff <= 24'd404577;
        419: data_ff <= -24'd259880;
        420: data_ff <= 24'd170580;
        421: data_ff <= -24'd111107;
        422: data_ff <= 24'd70571;
        423: data_ff <= -24'd43145;
        424: data_ff <= 24'd25092;
        425: data_ff <= -24'd13706;
        426: data_ff <= 24'd6923;
        427: data_ff <= -24'd3165;
        428: data_ff <= 24'd1268;
        429: data_ff <= -24'd417;
        430: data_ff <= 24'd93;
        431: data_ff <= -24'd7;
        432: data_ff <= 24'd1648472;
        433: data_ff <= -24'd711796;
        434: data_ff <= 24'd418965;
        435: data_ff <= -24'd268911;
        436: data_ff <= 24'd176416;
        437: data_ff <= -24'd114865;
        438: data_ff <= 24'd72938;
        439: data_ff <= -24'd44584;
        440: data_ff <= 24'd25926;
        441: data_ff <= -24'd14162;
        442: data_ff <= 24'd7154;
        443: data_ff <= -24'd3272;
        444: data_ff <= 24'd1311;
        445: data_ff <= -24'd432;
        446: data_ff <= 24'd97;
        447: data_ff <= -24'd7;
        448: data_ff <= 24'd1714652;
        449: data_ff <= -24'd737147;
        450: data_ff <= 24'd433276;
        451: data_ff <= -24'd277886;
        452: data_ff <= 24'd182215;
        453: data_ff <= -24'd118600;
        454: data_ff <= 24'd75291;
        455: data_ff <= -24'd46015;
        456: data_ff <= 24'd26756;
        457: data_ff <= -24'd14615;
        458: data_ff <= 24'd7384;
        459: data_ff <= -24'd3378;
        460: data_ff <= 24'd1354;
        461: data_ff <= -24'd447;
        462: data_ff <= 24'd101;
        463: data_ff <= -24'd8;
        464: data_ff <= 24'd1781204;
        465: data_ff <= -24'd762410;
        466: data_ff <= 24'd447503;
        467: data_ff <= -24'd286802;
        468: data_ff <= 24'd187973;
        469: data_ff <= -24'd122308;
        470: data_ff <= 24'd77628;
        471: data_ff <= -24'd47437;
        472: data_ff <= 24'd27581;
        473: data_ff <= -24'd15066;
        474: data_ff <= 24'd7613;
        475: data_ff <= -24'd3484;
        476: data_ff <= 24'd1398;
        477: data_ff <= -24'd462;
        478: data_ff <= 24'd104;
        479: data_ff <= -24'd8;
        480: data_ff <= 24'd1848116;
        481: data_ff <= -24'd787576;
        482: data_ff <= 24'd461642;
        483: data_ff <= -24'd295654;
        484: data_ff <= 24'd193689;
        485: data_ff <= -24'd125990;
        486: data_ff <= 24'd79949;
        487: data_ff <= -24'd48849;
        488: data_ff <= 24'd28401;
        489: data_ff <= -24'd15515;
        490: data_ff <= 24'd7842;
        491: data_ff <= -24'd3590;
        492: data_ff <= 24'd1441;
        493: data_ff <= -24'd476;
        494: data_ff <= 24'd108;
        495: data_ff <= -24'd8;
        496: data_ff <= 24'd1915376;
        497: data_ff <= -24'd812635;
        498: data_ff <= 24'd475687;
        499: data_ff <= -24'd304439;
        500: data_ff <= 24'd199360;
        501: data_ff <= -24'd129643;
        502: data_ff <= 24'd82252;
        503: data_ff <= -24'd50251;
        504: data_ff <= 24'd29216;
        505: data_ff <= -24'd15962;
        506: data_ff <= 24'd8069;
        507: data_ff <= -24'd3695;
        508: data_ff <= 24'd1484;
        509: data_ff <= -24'd491;
        510: data_ff <= 24'd112;
        511: data_ff <= -24'd9;
        512: data_ff <= 24'd1982970;
        513: data_ff <= -24'd837576;
        514: data_ff <= 24'd489630;
        515: data_ff <= -24'd313154;
        516: data_ff <= 24'd204984;
        517: data_ff <= -24'd133265;
        518: data_ff <= 24'd84536;
        519: data_ff <= -24'd51643;
        520: data_ff <= 24'd30025;
        521: data_ff <= -24'd16405;
        522: data_ff <= 24'd8295;
        523: data_ff <= -24'd3800;
        524: data_ff <= 24'd1527;
        525: data_ff <= -24'd506;
        526: data_ff <= 24'd116;
        527: data_ff <= -24'd9;
        528: data_ff <= 24'd2050886;
        529: data_ff <= -24'd862389;
        530: data_ff <= 24'd503467;
        531: data_ff <= -24'd321793;
        532: data_ff <= 24'd210557;
        533: data_ff <= -24'd136855;
        534: data_ff <= 24'd86801;
        535: data_ff <= -24'd53023;
        536: data_ff <= 24'd30828;
        537: data_ff <= -24'd16846;
        538: data_ff <= 24'd8519;
        539: data_ff <= -24'd3905;
        540: data_ff <= 24'd1570;
        541: data_ff <= -24'd521;
        542: data_ff <= 24'd120;
        543: data_ff <= -24'd9;
        544: data_ff <= 24'd2119110;
        545: data_ff <= -24'd887063;
        546: data_ff <= 24'd517191;
        547: data_ff <= -24'd330353;
        548: data_ff <= 24'd216079;
        549: data_ff <= -24'd140411;
        550: data_ff <= 24'd89045;
        551: data_ff <= -24'd54391;
        552: data_ff <= 24'd31624;
        553: data_ff <= -24'd17283;
        554: data_ff <= 24'd8742;
        555: data_ff <= -24'd4008;
        556: data_ff <= 24'd1613;
        557: data_ff <= -24'd536;
        558: data_ff <= 24'd123;
        559: data_ff <= -24'd10;
        560: data_ff <= 24'd2187630;
        561: data_ff <= -24'd911590;
        562: data_ff <= 24'd530796;
        563: data_ff <= -24'd338832;
        564: data_ff <= 24'd221545;
        565: data_ff <= -24'd143933;
        566: data_ff <= 24'd91267;
        567: data_ff <= -24'd55746;
        568: data_ff <= 24'd32414;
        569: data_ff <= -24'd17717;
        570: data_ff <= 24'd8964;
        571: data_ff <= -24'd4112;
        572: data_ff <= 24'd1656;
        573: data_ff <= -24'd551;
        574: data_ff <= 24'd127;
        575: data_ff <= -24'd10;
        576: data_ff <= 24'd2256431;
        577: data_ff <= -24'd935958;
        578: data_ff <= 24'd544277;
        579: data_ff <= -24'd347224;
        580: data_ff <= 24'd226954;
        581: data_ff <= -24'd147417;
        582: data_ff <= 24'd93467;
        583: data_ff <= -24'd57088;
        584: data_ff <= 24'd33196;
        585: data_ff <= -24'd18147;
        586: data_ff <= 24'd9184;
        587: data_ff <= -24'd4214;
        588: data_ff <= 24'd1698;
        589: data_ff <= -24'd566;
        590: data_ff <= 24'd131;
        591: data_ff <= -24'd10;
        592: data_ff <= 24'd2325500;
        593: data_ff <= -24'd960157;
        594: data_ff <= 24'd557627;
        595: data_ff <= -24'd355527;
        596: data_ff <= 24'd232303;
        597: data_ff <= -24'd150863;
        598: data_ff <= 24'd95642;
        599: data_ff <= -24'd58416;
        600: data_ff <= 24'd33970;
        601: data_ff <= -24'd18573;
        602: data_ff <= 24'd9402;
        603: data_ff <= -24'd4316;
        604: data_ff <= 24'd1741;
        605: data_ff <= -24'd581;
        606: data_ff <= 24'd135;
        607: data_ff <= -24'd11;
        608: data_ff <= 24'd2394824;
        609: data_ff <= -24'd984176;
        610: data_ff <= 24'd570841;
        611: data_ff <= -24'd363735;
        612: data_ff <= 24'd237590;
        613: data_ff <= -24'd154269;
        614: data_ff <= 24'd97794;
        615: data_ff <= -24'd59730;
        616: data_ff <= 24'd34737;
        617: data_ff <= -24'd18995;
        618: data_ff <= 24'd9619;
        619: data_ff <= -24'd4418;
        620: data_ff <= 24'd1783;
        621: data_ff <= -24'd595;
        622: data_ff <= 24'd139;
        623: data_ff <= -24'd11;
        624: data_ff <= 24'd2464388;
        625: data_ff <= -24'd1008006;
        626: data_ff <= 24'd583912;
        627: data_ff <= -24'd371847;
        628: data_ff <= 24'd242812;
        629: data_ff <= -24'd157633;
        630: data_ff <= 24'd99919;
        631: data_ff <= -24'd61029;
        632: data_ff <= 24'd35495;
        633: data_ff <= -24'd19413;
        634: data_ff <= 24'd9833;
        635: data_ff <= -24'd4518;
        636: data_ff <= 24'd1825;
        637: data_ff <= -24'd610;
        638: data_ff <= 24'd143;
        639: data_ff <= -24'd12;
        640: data_ff <= 24'd2534180;
        641: data_ff <= -24'd1031637;
        642: data_ff <= 24'd596835;
        643: data_ff <= -24'd379858;
        644: data_ff <= 24'd247968;
        645: data_ff <= -24'd160954;
        646: data_ff <= 24'd102018;
        647: data_ff <= -24'd62311;
        648: data_ff <= 24'd36244;
        649: data_ff <= -24'd19827;
        650: data_ff <= 24'd10045;
        651: data_ff <= -24'd4618;
        652: data_ff <= 24'd1866;
        653: data_ff <= -24'd625;
        654: data_ff <= 24'd147;
        655: data_ff <= -24'd12;
        656: data_ff <= 24'd2604185;
        657: data_ff <= -24'd1055057;
        658: data_ff <= 24'd609604;
        659: data_ff <= -24'd387764;
        660: data_ff <= 24'd253054;
        661: data_ff <= -24'd164230;
        662: data_ff <= 24'd104088;
        663: data_ff <= -24'd63578;
        664: data_ff <= 24'd36985;
        665: data_ff <= -24'd20235;
        666: data_ff <= 24'd10256;
        667: data_ff <= -24'd4717;
        668: data_ff <= 24'd1907;
        669: data_ff <= -24'd639;
        670: data_ff <= 24'd151;
        671: data_ff <= -24'd13;
        672: data_ff <= 24'd2674389;
        673: data_ff <= -24'd1078257;
        674: data_ff <= 24'd622212;
        675: data_ff <= -24'd395561;
        676: data_ff <= 24'd258068;
        677: data_ff <= -24'd167461;
        678: data_ff <= 24'd106131;
        679: data_ff <= -24'd64827;
        680: data_ff <= 24'd37716;
        681: data_ff <= -24'd20639;
        682: data_ff <= 24'd10463;
        683: data_ff <= -24'd4814;
        684: data_ff <= 24'd1948;
        685: data_ff <= -24'd654;
        686: data_ff <= 24'd155;
        687: data_ff <= -24'd13;
        688: data_ff <= 24'd2744777;
        689: data_ff <= -24'd1101225;
        690: data_ff <= 24'd634655;
        691: data_ff <= -24'd403247;
        692: data_ff <= 24'd263008;
        693: data_ff <= -24'd170643;
        694: data_ff <= 24'd108143;
        695: data_ff <= -24'd66059;
        696: data_ff <= 24'd38437;
        697: data_ff <= -24'd21038;
        698: data_ff <= 24'd10669;
        699: data_ff <= -24'd4911;
        700: data_ff <= 24'd1989;
        701: data_ff <= -24'd668;
        702: data_ff <= 24'd158;
        703: data_ff <= -24'd13;
        704: data_ff <= 24'd2815337;
        705: data_ff <= -24'd1123953;
        706: data_ff <= 24'd646927;
        707: data_ff <= -24'd410817;
        708: data_ff <= 24'd267872;
        709: data_ff <= -24'd173776;
        710: data_ff <= 24'd110125;
        711: data_ff <= -24'd67272;
        712: data_ff <= 24'd39147;
        713: data_ff <= -24'd21432;
        714: data_ff <= 24'd10872;
        715: data_ff <= -24'd5007;
        716: data_ff <= 24'd2029;
        717: data_ff <= -24'd683;
        718: data_ff <= 24'd162;
        719: data_ff <= -24'd14;
        720: data_ff <= 24'd2886052;
        721: data_ff <= -24'd1146429;
        722: data_ff <= 24'd659021;
        723: data_ff <= -24'd418268;
        724: data_ff <= 24'd272657;
        725: data_ff <= -24'd176858;
        726: data_ff <= 24'd112075;
        727: data_ff <= -24'd68467;
        728: data_ff <= 24'd39848;
        729: data_ff <= -24'd21820;
        730: data_ff <= 24'd11072;
        731: data_ff <= -24'd5102;
        732: data_ff <= 24'd2069;
        733: data_ff <= -24'd697;
        734: data_ff <= 24'd166;
        735: data_ff <= -24'd14;
        736: data_ff <= 24'd2956910;
        737: data_ff <= -24'd1168642;
        738: data_ff <= 24'd670931;
        739: data_ff <= -24'd425597;
        740: data_ff <= 24'd277361;
        741: data_ff <= -24'd179888;
        742: data_ff <= 24'd113993;
        743: data_ff <= -24'd69643;
        744: data_ff <= 24'd40537;
        745: data_ff <= -24'd22202;
        746: data_ff <= 24'd11270;
        747: data_ff <= -24'd5195;
        748: data_ff <= 24'd2109;
        749: data_ff <= -24'd711;
        750: data_ff <= 24'd170;
        751: data_ff <= -24'd15;
        752: data_ff <= 24'd3027895;
        753: data_ff <= -24'd1190584;
        754: data_ff <= 24'd682653;
        755: data_ff <= -24'd432799;
        756: data_ff <= 24'd281982;
        757: data_ff <= -24'd182864;
        758: data_ff <= 24'd115877;
        759: data_ff <= -24'd70798;
        760: data_ff <= 24'd41215;
        761: data_ff <= -24'd22578;
        762: data_ff <= 24'd11465;
        763: data_ff <= -24'd5288;
        764: data_ff <= 24'd2148;
        765: data_ff <= -24'd726;
        766: data_ff <= 24'd174;
        767: data_ff <= -24'd15;
        768: data_ff <= 24'd3098993;
        769: data_ff <= -24'd1212243;
        770: data_ff <= 24'd694181;
        771: data_ff <= -24'd439872;
        772: data_ff <= 24'd286517;
        773: data_ff <= -24'd185785;
        774: data_ff <= 24'd117726;
        775: data_ff <= -24'd71932;
        776: data_ff <= 24'd41882;
        777: data_ff <= -24'd22949;
        778: data_ff <= 24'd11657;
        779: data_ff <= -24'd5379;
        780: data_ff <= 24'd2187;
        781: data_ff <= -24'd740;
        782: data_ff <= 24'd178;
        783: data_ff <= -24'd16;
        784: data_ff <= 24'd3170189;
        785: data_ff <= -24'd1233609;
        786: data_ff <= 24'd705508;
        787: data_ff <= -24'd446811;
        788: data_ff <= 24'd290964;
        789: data_ff <= -24'd188649;
        790: data_ff <= 24'd119540;
        791: data_ff <= -24'd73046;
        792: data_ff <= 24'd42536;
        793: data_ff <= -24'd23313;
        794: data_ff <= 24'd11846;
        795: data_ff <= -24'd5469;
        796: data_ff <= 24'd2225;
        797: data_ff <= -24'd753;
        798: data_ff <= 24'd182;
        799: data_ff <= -24'd16;
        800: data_ff <= 24'd3241469;
        801: data_ff <= -24'd1254672;
        802: data_ff <= 24'd716630;
        803: data_ff <= -24'd453614;
        804: data_ff <= 24'd295321;
        805: data_ff <= -24'd191455;
        806: data_ff <= 24'd121317;
        807: data_ff <= -24'd74138;
        808: data_ff <= 24'd43179;
        809: data_ff <= -24'd23670;
        810: data_ff <= 24'd12032;
        811: data_ff <= -24'd5557;
        812: data_ff <= 24'd2262;
        813: data_ff <= -24'd767;
        814: data_ff <= 24'd186;
        815: data_ff <= -24'd17;
        816: data_ff <= 24'd3312817;
        817: data_ff <= -24'd1275421;
        818: data_ff <= 24'd727540;
        819: data_ff <= -24'd460276;
        820: data_ff <= 24'd299585;
        821: data_ff <= -24'd194201;
        822: data_ff <= 24'd123058;
        823: data_ff <= -24'd75207;
        824: data_ff <= 24'd43808;
        825: data_ff <= -24'd24021;
        826: data_ff <= 24'd12214;
        827: data_ff <= -24'd5645;
        828: data_ff <= 24'd2300;
        829: data_ff <= -24'd781;
        830: data_ff <= 24'd190;
        831: data_ff <= -24'd17;
        832: data_ff <= 24'd3384219;
        833: data_ff <= -24'd1295847;
        834: data_ff <= 24'd738234;
        835: data_ff <= -24'd466796;
        836: data_ff <= 24'd303756;
        837: data_ff <= -24'd196886;
        838: data_ff <= 24'd124760;
        839: data_ff <= -24'd76253;
        840: data_ff <= 24'd44425;
        841: data_ff <= -24'd24365;
        842: data_ff <= 24'd12394;
        843: data_ff <= -24'd5730;
        844: data_ff <= 24'd2336;
        845: data_ff <= -24'd794;
        846: data_ff <= 24'd193;
        847: data_ff <= -24'd18;
        848: data_ff <= 24'd3455661;
        849: data_ff <= -24'd1315938;
        850: data_ff <= 24'd748705;
        851: data_ff <= -24'd473168;
        852: data_ff <= 24'd307829;
        853: data_ff <= -24'd199509;
        854: data_ff <= 24'd126422;
        855: data_ff <= -24'd77276;
        856: data_ff <= 24'd45028;
        857: data_ff <= -24'd24702;
        858: data_ff <= 24'd12569;
        859: data_ff <= -24'd5815;
        860: data_ff <= 24'd2372;
        861: data_ff <= -24'd807;
        862: data_ff <= 24'd197;
        863: data_ff <= -24'd18;
        864: data_ff <= 24'd3527126;
        865: data_ff <= -24'd1335686;
        866: data_ff <= 24'd758949;
        867: data_ff <= -24'd479391;
        868: data_ff <= 24'd311804;
        869: data_ff <= -24'd202067;
        870: data_ff <= 24'd128045;
        871: data_ff <= -24'd78275;
        872: data_ff <= 24'd45617;
        873: data_ff <= -24'd25032;
        874: data_ff <= 24'd12742;
        875: data_ff <= -24'd5897;
        876: data_ff <= 24'd2408;
        877: data_ff <= -24'd821;
        878: data_ff <= 24'd201;
        879: data_ff <= -24'd19;
        880: data_ff <= 24'd3598600;
        881: data_ff <= -24'd1355079;
        882: data_ff <= 24'd768960;
        883: data_ff <= -24'd485460;
        884: data_ff <= 24'd315679;
        885: data_ff <= -24'd204561;
        886: data_ff <= 24'd129627;
        887: data_ff <= -24'd79249;
        888: data_ff <= 24'd46193;
        889: data_ff <= -24'd25354;
        890: data_ff <= 24'd12910;
        891: data_ff <= -24'd5978;
        892: data_ff <= 24'd2443;
        893: data_ff <= -24'd834;
        894: data_ff <= 24'd205;
        895: data_ff <= -24'd19;
        896: data_ff <= 24'd3670068;
        897: data_ff <= -24'd1374108;
        898: data_ff <= 24'd778733;
        899: data_ff <= -24'd491373;
        900: data_ff <= 24'd319450;
        901: data_ff <= -24'd206988;
        902: data_ff <= 24'd131167;
        903: data_ff <= -24'd80198;
        904: data_ff <= 24'd46754;
        905: data_ff <= -24'd25668;
        906: data_ff <= 24'd13075;
        907: data_ff <= -24'd6058;
        908: data_ff <= 24'd2477;
        909: data_ff <= -24'd846;
        910: data_ff <= 24'd209;
        911: data_ff <= -24'd20;
        912: data_ff <= 24'd3741515;
        913: data_ff <= -24'd1392762;
        914: data_ff <= 24'd788262;
        915: data_ff <= -24'd497126;
        916: data_ff <= 24'd323116;
        917: data_ff <= -24'd209347;
        918: data_ff <= 24'd132664;
        919: data_ff <= -24'd81122;
        920: data_ff <= 24'd47300;
        921: data_ff <= -24'd25975;
        922: data_ff <= 24'd13236;
        923: data_ff <= -24'd6135;
        924: data_ff <= 24'd2511;
        925: data_ff <= -24'd859;
        926: data_ff <= 24'd212;
        927: data_ff <= -24'd21;
        928: data_ff <= 24'd3812926;
        929: data_ff <= -24'd1411032;
        930: data_ff <= 24'd797543;
        931: data_ff <= -24'd502717;
        932: data_ff <= 24'd326676;
        933: data_ff <= -24'd211637;
        934: data_ff <= 24'd134118;
        935: data_ff <= -24'd82019;
        936: data_ff <= 24'd47831;
        937: data_ff <= -24'd26273;
        938: data_ff <= 24'd13393;
        939: data_ff <= -24'd6211;
        940: data_ff <= 24'd2544;
        941: data_ff <= -24'd871;
        942: data_ff <= 24'd216;
        943: data_ff <= -24'd21;
        944: data_ff <= 24'd3884285;
        945: data_ff <= -24'd1428907;
        946: data_ff <= 24'd806570;
        947: data_ff <= -24'd508142;
        948: data_ff <= 24'd330126;
        949: data_ff <= -24'd213856;
        950: data_ff <= 24'd135528;
        951: data_ff <= -24'd82889;
        952: data_ff <= 24'd48347;
        953: data_ff <= -24'd26563;
        954: data_ff <= 24'd13546;
        955: data_ff <= -24'd6285;
        956: data_ff <= 24'd2576;
        957: data_ff <= -24'd883;
        958: data_ff <= 24'd220;
        959: data_ff <= -24'd22;
        960: data_ff <= 24'd3955577;
        961: data_ff <= -24'd1446378;
        962: data_ff <= 24'd815339;
        963: data_ff <= -24'd513398;
        964: data_ff <= 24'd333466;
        965: data_ff <= -24'd216004;
        966: data_ff <= 24'd136892;
        967: data_ff <= -24'd83732;
        968: data_ff <= 24'd48848;
        969: data_ff <= -24'd26845;
        970: data_ff <= 24'd13694;
        971: data_ff <= -24'd6358;
        972: data_ff <= 24'd2608;
        973: data_ff <= -24'd895;
        974: data_ff <= 24'd223;
        975: data_ff <= -24'd22;
        976: data_ff <= 24'd4026788;
        977: data_ff <= -24'd1463435;
        978: data_ff <= 24'd823843;
        979: data_ff <= -24'd518482;
        980: data_ff <= 24'd336693;
        981: data_ff <= -24'd218079;
        982: data_ff <= 24'd138210;
        983: data_ff <= -24'd84547;
        984: data_ff <= 24'd49332;
        985: data_ff <= -24'd27119;
        986: data_ff <= 24'd13839;
        987: data_ff <= -24'd6428;
        988: data_ff <= 24'd2638;
        989: data_ff <= -24'd907;
        990: data_ff <= 24'd227;
        991: data_ff <= -24'd23;
        992: data_ff <= 24'd4097901;
        993: data_ff <= -24'd1480067;
        994: data_ff <= 24'd832079;
        995: data_ff <= -24'd523391;
        996: data_ff <= 24'd339805;
        997: data_ff <= -24'd220079;
        998: data_ff <= 24'd139482;
        999: data_ff <= -24'd85334;
        1000: data_ff <= 24'd49800;
        1001: data_ff <= -24'd27383;
        1002: data_ff <= 24'd13979;
        1003: data_ff <= -24'd6496;
        1004: data_ff <= 24'd2669;
        1005: data_ff <= -24'd919;
        1006: data_ff <= 24'd230;
        1007: data_ff <= -24'd23;
        1008: data_ff <= 24'd4168902;
        1009: data_ff <= -24'd1496266;
        1010: data_ff <= 24'd840042;
        1011: data_ff <= -24'd528123;
        1012: data_ff <= 24'd342801;
        1013: data_ff <= -24'd222004;
        1014: data_ff <= 24'd140706;
        1015: data_ff <= -24'd86092;
        1016: data_ff <= 24'd50251;
        1017: data_ff <= -24'd27639;
        1018: data_ff <= 24'd14115;
        1019: data_ff <= -24'd6563;
        1020: data_ff <= 24'd2698;
        1021: data_ff <= -24'd930;
        1022: data_ff <= 24'd234;
        1023: data_ff <= -24'd24;
        1024: data_ff <= 24'd4239775;
        1025: data_ff <= -24'd1512022;
        1026: data_ff <= 24'd847726;
        1027: data_ff <= -24'd532674;
        1028: data_ff <= 24'd345679;
        1029: data_ff <= -24'd223852;
        1030: data_ff <= 24'd141882;
        1031: data_ff <= -24'd86821;
        1032: data_ff <= 24'd50686;
        1033: data_ff <= -24'd27885;
        1034: data_ff <= 24'd14246;
        1035: data_ff <= -24'd6627;
        1036: data_ff <= 24'd2726;
        1037: data_ff <= -24'd941;
        1038: data_ff <= 24'd237;
        1039: data_ff <= -24'd24;
        1040: data_ff <= 24'd4310505;
        1041: data_ff <= -24'd1527324;
        1042: data_ff <= 24'd855127;
        1043: data_ff <= -24'd537042;
        1044: data_ff <= 24'd348437;
        1045: data_ff <= -24'd225623;
        1046: data_ff <= 24'd143009;
        1047: data_ff <= -24'd87520;
        1048: data_ff <= 24'd51103;
        1049: data_ff <= -24'd28122;
        1050: data_ff <= 24'd14372;
        1051: data_ff <= -24'd6690;
        1052: data_ff <= 24'd2754;
        1053: data_ff <= -24'd951;
        1054: data_ff <= 24'd241;
        1055: data_ff <= -24'd25;
        1056: data_ff <= 24'd4381077;
        1057: data_ff <= -24'd1542164;
        1058: data_ff <= 24'd862241;
        1059: data_ff <= -24'd541224;
        1060: data_ff <= 24'd351073;
        1061: data_ff <= -24'd227315;
        1062: data_ff <= 24'd144085;
        1063: data_ff <= -24'd88188;
        1064: data_ff <= 24'd51503;
        1065: data_ff <= -24'd28350;
        1066: data_ff <= 24'd14494;
        1067: data_ff <= -24'd6750;
        1068: data_ff <= 24'd2781;
        1069: data_ff <= -24'd962;
        1070: data_ff <= 24'd244;
        1071: data_ff <= -24'd26;
        1072: data_ff <= 24'd4451475;
        1073: data_ff <= -24'd1556531;
        1074: data_ff <= 24'd869063;
        1075: data_ff <= -24'd545218;
        1076: data_ff <= 24'd353585;
        1077: data_ff <= -24'd228926;
        1078: data_ff <= 24'd145112;
        1079: data_ff <= -24'd88826;
        1080: data_ff <= 24'd51885;
        1081: data_ff <= -24'd28568;
        1082: data_ff <= 24'd14611;
        1083: data_ff <= -24'd6808;
        1084: data_ff <= 24'd2807;
        1085: data_ff <= -24'd972;
        1086: data_ff <= 24'd247;
        1087: data_ff <= -24'd26;
        1088: data_ff <= 24'd4521684;
        1089: data_ff <= -24'd1570418;
        1090: data_ff <= 24'd875588;
        1091: data_ff <= -24'd549020;
        1092: data_ff <= 24'd355973;
        1093: data_ff <= -24'd230457;
        1094: data_ff <= 24'd146087;
        1095: data_ff <= -24'd89433;
        1096: data_ff <= 24'd52250;
        1097: data_ff <= -24'd28776;
        1098: data_ff <= 24'd14723;
        1099: data_ff <= -24'd6863;
        1100: data_ff <= 24'd2832;
        1101: data_ff <= -24'd982;
        1102: data_ff <= 24'd250;
        1103: data_ff <= -24'd27;
        1104: data_ff <= 24'd4591688;
        1105: data_ff <= -24'd1583813;
        1106: data_ff <= 24'd881812;
        1107: data_ff <= -24'd552629;
        1108: data_ff <= 24'd358233;
        1109: data_ff <= -24'd231905;
        1110: data_ff <= 24'd147010;
        1111: data_ff <= -24'd90008;
        1112: data_ff <= 24'd52595;
        1113: data_ff <= -24'd28974;
        1114: data_ff <= 24'd14830;
        1115: data_ff <= -24'd6917;
        1116: data_ff <= 24'd2856;
        1117: data_ff <= -24'd992;
        1118: data_ff <= 24'd253;
        1119: data_ff <= -24'd27;
        1120: data_ff <= 24'd4661473;
        1121: data_ff <= -24'd1596708;
        1122: data_ff <= 24'd887731;
        1123: data_ff <= -24'd556041;
        1124: data_ff <= 24'd360366;
        1125: data_ff <= -24'd233271;
        1126: data_ff <= 24'd147880;
        1127: data_ff <= -24'd90551;
        1128: data_ff <= 24'd52923;
        1129: data_ff <= -24'd29162;
        1130: data_ff <= 24'd14931;
        1131: data_ff <= -24'd6968;
        1132: data_ff <= 24'd2879;
        1133: data_ff <= -24'd1001;
        1134: data_ff <= 24'd256;
        1135: data_ff <= -24'd28;
        1136: data_ff <= 24'd4731023;
        1137: data_ff <= -24'd1609095;
        1138: data_ff <= 24'd893341;
        1139: data_ff <= -24'd559255;
        1140: data_ff <= 24'd362368;
        1141: data_ff <= -24'd234552;
        1142: data_ff <= 24'd148698;
        1143: data_ff <= -24'd91062;
        1144: data_ff <= 24'd53231;
        1145: data_ff <= -24'd29340;
        1146: data_ff <= 24'd15028;
        1147: data_ff <= -24'd7016;
        1148: data_ff <= 24'd2902;
        1149: data_ff <= -24'd1010;
        1150: data_ff <= 24'd259;
        1151: data_ff <= -24'd29;
        1152: data_ff <= 24'd4800323;
        1153: data_ff <= -24'd1620963;
        1154: data_ff <= 24'd898637;
        1155: data_ff <= -24'd562268;
        1156: data_ff <= 24'd364240;
        1157: data_ff <= -24'd235748;
        1158: data_ff <= 24'd149461;
        1159: data_ff <= -24'd91540;
        1160: data_ff <= 24'd53520;
        1161: data_ff <= -24'd29507;
        1162: data_ff <= 24'd15119;
        1163: data_ff <= -24'd7063;
        1164: data_ff <= 24'd2923;
        1165: data_ff <= -24'd1018;
        1166: data_ff <= 24'd262;
        1167: data_ff <= -24'd29;
        1168: data_ff <= 24'd4869357;
        1169: data_ff <= -24'd1632304;
        1170: data_ff <= 24'd903615;
        1171: data_ff <= -24'd565077;
        1172: data_ff <= 24'd365978;
        1173: data_ff <= -24'd236858;
        1174: data_ff <= 24'd150170;
        1175: data_ff <= -24'd91984;
        1176: data_ff <= 24'd53790;
        1177: data_ff <= -24'd29664;
        1178: data_ff <= 24'd15205;
        1179: data_ff <= -24'd7106;
        1180: data_ff <= 24'd2943;
        1181: data_ff <= -24'd1027;
        1182: data_ff <= 24'd265;
        1183: data_ff <= -24'd30;
        1184: data_ff <= 24'd4938111;
        1185: data_ff <= -24'd1643109;
        1186: data_ff <= 24'd908272;
        1187: data_ff <= -24'd567682;
        1188: data_ff <= 24'd367583;
        1189: data_ff <= -24'd237881;
        1190: data_ff <= 24'd150824;
        1191: data_ff <= -24'd92395;
        1192: data_ff <= 24'd54040;
        1193: data_ff <= -24'd29810;
        1194: data_ff <= 24'd15286;
        1195: data_ff <= -24'd7148;
        1196: data_ff <= 24'd2962;
        1197: data_ff <= -24'd1035;
        1198: data_ff <= 24'd268;
        1199: data_ff <= -24'd30;
        1200: data_ff <= 24'd5006569;
        1201: data_ff <= -24'd1653370;
        1202: data_ff <= 24'd912604;
        1203: data_ff <= -24'd570078;
        1204: data_ff <= 24'd369052;
        1205: data_ff <= -24'd238815;
        1206: data_ff <= 24'd151422;
        1207: data_ff <= -24'd92772;
        1208: data_ff <= 24'd54271;
        1209: data_ff <= -24'd29945;
        1210: data_ff <= 24'd15361;
        1211: data_ff <= -24'd7186;
        1212: data_ff <= 24'd2981;
        1213: data_ff <= -24'd1042;
        1214: data_ff <= 24'd271;
        1215: data_ff <= -24'd31;
        1216: data_ff <= 24'd5074717;
        1217: data_ff <= -24'd1663077;
        1218: data_ff <= 24'd916607;
        1219: data_ff <= -24'd572265;
        1220: data_ff <= 24'd370384;
        1221: data_ff <= -24'd239662;
        1222: data_ff <= 24'd151963;
        1223: data_ff <= -24'd93114;
        1224: data_ff <= 24'd54481;
        1225: data_ff <= -24'd30069;
        1226: data_ff <= 24'd15430;
        1227: data_ff <= -24'd7223;
        1228: data_ff <= 24'd2998;
        1229: data_ff <= -24'd1050;
        1230: data_ff <= 24'd273;
        1231: data_ff <= -24'd31;
        1232: data_ff <= 24'd5142538;
        1233: data_ff <= -24'd1672222;
        1234: data_ff <= 24'd920277;
        1235: data_ff <= -24'd574240;
        1236: data_ff <= 24'd371578;
        1237: data_ff <= -24'd240418;
        1238: data_ff <= 24'd152448;
        1239: data_ff <= -24'd93422;
        1240: data_ff <= 24'd54671;
        1241: data_ff <= -24'd30182;
        1242: data_ff <= 24'd15494;
        1243: data_ff <= -24'd7256;
        1244: data_ff <= 24'd3014;
        1245: data_ff <= -24'd1056;
        1246: data_ff <= 24'd276;
        1247: data_ff <= -24'd32;
        1248: data_ff <= 24'd5210018;
        1249: data_ff <= -24'd1680797;
        1250: data_ff <= 24'd923611;
        1251: data_ff <= -24'd576001;
        1252: data_ff <= 24'd372633;
        1253: data_ff <= -24'd241085;
        1254: data_ff <= 24'd152876;
        1255: data_ff <= -24'd93694;
        1256: data_ff <= 24'd54841;
        1257: data_ff <= -24'd30284;
        1258: data_ff <= 24'd15552;
        1259: data_ff <= -24'd7287;
        1260: data_ff <= 24'd3029;
        1261: data_ff <= -24'd1063;
        1262: data_ff <= 24'd278;
        1263: data_ff <= -24'd33;
        1264: data_ff <= 24'd5277142;
        1265: data_ff <= -24'd1688793;
        1266: data_ff <= 24'd926606;
        1267: data_ff <= -24'd577547;
        1268: data_ff <= 24'd373547;
        1269: data_ff <= -24'd241660;
        1270: data_ff <= 24'd153246;
        1271: data_ff <= -24'd93931;
        1272: data_ff <= 24'd54990;
        1273: data_ff <= -24'd30374;
        1274: data_ff <= 24'd15604;
        1275: data_ff <= -24'd7315;
        1276: data_ff <= 24'd3043;
        1277: data_ff <= -24'd1069;
        1278: data_ff <= 24'd280;
        1279: data_ff <= -24'd33;
        1280: data_ff <= 24'd5343894;
        1281: data_ff <= -24'd1696203;
        1282: data_ff <= 24'd929257;
        1283: data_ff <= -24'd578875;
        1284: data_ff <= 24'd374320;
        1285: data_ff <= -24'd242143;
        1286: data_ff <= 24'd153557;
        1287: data_ff <= -24'd94133;
        1288: data_ff <= 24'd55118;
        1289: data_ff <= -24'd30453;
        1290: data_ff <= 24'd15650;
        1291: data_ff <= -24'd7340;
        1292: data_ff <= 24'd3056;
        1293: data_ff <= -24'd1075;
        1294: data_ff <= 24'd283;
        1295: data_ff <= -24'd34;
        1296: data_ff <= 24'd5410261;
        1297: data_ff <= -24'd1703018;
        1298: data_ff <= 24'd931562;
        1299: data_ff <= -24'd579984;
        1300: data_ff <= 24'd374951;
        1301: data_ff <= -24'd242534;
        1302: data_ff <= 24'd153810;
        1303: data_ff <= -24'd94298;
        1304: data_ff <= 24'd55224;
        1305: data_ff <= -24'd30520;
        1306: data_ff <= 24'd15690;
        1307: data_ff <= -24'd7363;
        1308: data_ff <= 24'd3067;
        1309: data_ff <= -24'd1080;
        1310: data_ff <= 24'd285;
        1311: data_ff <= -24'd34;
        1312: data_ff <= 24'd5476227;
        1313: data_ff <= -24'd1709230;
        1314: data_ff <= 24'd933519;
        1315: data_ff <= -24'd580873;
        1316: data_ff <= 24'd375437;
        1317: data_ff <= -24'd242832;
        1318: data_ff <= 24'd154003;
        1319: data_ff <= -24'd94427;
        1320: data_ff <= 24'd55310;
        1321: data_ff <= -24'd30575;
        1322: data_ff <= 24'd15724;
        1323: data_ff <= -24'd7383;
        1324: data_ff <= 24'd3078;
        1325: data_ff <= -24'd1085;
        1326: data_ff <= 24'd287;
        1327: data_ff <= -24'd35;
        1328: data_ff <= 24'd5541777;
        1329: data_ff <= -24'd1714832;
        1330: data_ff <= 24'd935122;
        1331: data_ff <= -24'd581539;
        1332: data_ff <= 24'd375779;
        1333: data_ff <= -24'd243035;
        1334: data_ff <= 24'd154137;
        1335: data_ff <= -24'd94519;
        1336: data_ff <= 24'd55374;
        1337: data_ff <= -24'd30618;
        1338: data_ff <= 24'd15752;
        1339: data_ff <= -24'd7399;
        1340: data_ff <= 24'd3087;
        1341: data_ff <= -24'd1090;
        1342: data_ff <= 24'd289;
        1343: data_ff <= -24'd35;
        1344: data_ff <= 24'd5606897;
        1345: data_ff <= -24'd1719815;
        1346: data_ff <= 24'd936371;
        1347: data_ff <= -24'd581982;
        1348: data_ff <= 24'd375976;
        1349: data_ff <= -24'd243145;
        1350: data_ff <= 24'd154210;
        1351: data_ff <= -24'd94574;
        1352: data_ff <= 24'd55416;
        1353: data_ff <= -24'd30650;
        1354: data_ff <= 24'd15774;
        1355: data_ff <= -24'd7413;
        1356: data_ff <= 24'd3095;
        1357: data_ff <= -24'd1094;
        1358: data_ff <= 24'd290;
        1359: data_ff <= -24'd36;
        1360: data_ff <= 24'd5671572;
        1361: data_ff <= -24'd1724172;
        1362: data_ff <= 24'd937262;
        1363: data_ff <= -24'd582199;
        1364: data_ff <= 24'd376026;
        1365: data_ff <= -24'd243159;
        1366: data_ff <= 24'd154223;
        1367: data_ff <= -24'd94592;
        1368: data_ff <= 24'd55437;
        1369: data_ff <= -24'd30669;
        1370: data_ff <= 24'd15790;
        1371: data_ff <= -24'd7424;
        1372: data_ff <= 24'd3102;
        1373: data_ff <= -24'd1097;
        1374: data_ff <= 24'd292;
        1375: data_ff <= -24'd36;
        1376: data_ff <= 24'd5735787;
        1377: data_ff <= -24'd1727896;
        1378: data_ff <= 24'd937792;
        1379: data_ff <= -24'd582189;
        1380: data_ff <= 24'd375930;
        1381: data_ff <= -24'd243077;
        1382: data_ff <= 24'd154176;
        1383: data_ff <= -24'd94572;
        1384: data_ff <= 24'd55435;
        1385: data_ff <= -24'd30676;
        1386: data_ff <= 24'd15799;
        1387: data_ff <= -24'd7432;
        1388: data_ff <= 24'd3107;
        1389: data_ff <= -24'd1100;
        1390: data_ff <= 24'd294;
        1391: data_ff <= -24'd37;
        1392: data_ff <= 24'd5799529;
        1393: data_ff <= -24'd1730980;
        1394: data_ff <= 24'd937959;
        1395: data_ff <= -24'd581952;
        1396: data_ff <= 24'd375685;
        1397: data_ff <= -24'd242900;
        1398: data_ff <= 24'd154067;
        1399: data_ff <= -24'd94515;
        1400: data_ff <= 24'd55411;
        1401: data_ff <= -24'd30671;
        1402: data_ff <= 24'd15802;
        1403: data_ff <= -24'd7437;
        1404: data_ff <= 24'd3112;
        1405: data_ff <= -24'd1103;
        1406: data_ff <= 24'd295;
        1407: data_ff <= -24'd37;
        1408: data_ff <= 24'd5862781;
        1409: data_ff <= -24'd1733415;
        1410: data_ff <= 24'd937761;
        1411: data_ff <= -24'd581486;
        1412: data_ff <= 24'd375291;
        1413: data_ff <= -24'd242626;
        1414: data_ff <= 24'd153897;
        1415: data_ff <= -24'd94420;
        1416: data_ff <= 24'd55365;
        1417: data_ff <= -24'd30653;
        1418: data_ff <= 24'd15798;
        1419: data_ff <= -24'd7439;
        1420: data_ff <= 24'd3115;
        1421: data_ff <= -24'd1106;
        1422: data_ff <= 24'd296;
        1423: data_ff <= -24'd38;
        1424: data_ff <= 24'd5925531;
        1425: data_ff <= -24'd1735196;
        1426: data_ff <= 24'd937195;
        1427: data_ff <= -24'd580789;
        1428: data_ff <= 24'd374749;
        1429: data_ff <= -24'd242256;
        1430: data_ff <= 24'd153665;
        1431: data_ff <= -24'd94287;
        1432: data_ff <= 24'd55297;
        1433: data_ff <= -24'd30623;
        1434: data_ff <= 24'd15788;
        1435: data_ff <= -24'd7438;
        1436: data_ff <= 24'd3116;
        1437: data_ff <= -24'd1107;
        1438: data_ff <= 24'd297;
        1439: data_ff <= -24'd38;
        1440: data_ff <= 24'd5987764;
        1441: data_ff <= -24'd1736316;
        1442: data_ff <= 24'd936258;
        1443: data_ff <= -24'd579862;
        1444: data_ff <= 24'd374056;
        1445: data_ff <= -24'd241787;
        1446: data_ff <= 24'd153371;
        1447: data_ff <= -24'd94116;
        1448: data_ff <= 24'd55206;
        1449: data_ff <= -24'd30580;
        1450: data_ff <= 24'd15771;
        1451: data_ff <= -24'd7434;
        1452: data_ff <= 24'd3117;
        1453: data_ff <= -24'd1109;
        1454: data_ff <= 24'd299;
        1455: data_ff <= -24'd39;
        1456: data_ff <= 24'd6049466;
        1457: data_ff <= -24'd1736767;
        1458: data_ff <= 24'd934950;
        1459: data_ff <= -24'd578702;
        1460: data_ff <= 24'd373213;
        1461: data_ff <= -24'd241222;
        1462: data_ff <= 24'd153014;
        1463: data_ff <= -24'd93906;
        1464: data_ff <= 24'd55092;
        1465: data_ff <= -24'd30524;
        1466: data_ff <= 24'd15748;
        1467: data_ff <= -24'd7427;
        1468: data_ff <= 24'd3116;
        1469: data_ff <= -24'd1110;
        1470: data_ff <= 24'd299;
        1471: data_ff <= -24'd39;
        1472: data_ff <= 24'd6110623;
        1473: data_ff <= -24'd1736543;
        1474: data_ff <= 24'd933268;
        1475: data_ff <= -24'd577309;
        1476: data_ff <= 24'd372219;
        1477: data_ff <= -24'd240558;
        1478: data_ff <= 24'd152595;
        1479: data_ff <= -24'd93658;
        1480: data_ff <= 24'd54955;
        1481: data_ff <= -24'd30456;
        1482: data_ff <= 24'd15718;
        1483: data_ff <= -24'd7416;
        1484: data_ff <= 24'd3114;
        1485: data_ff <= -24'd1110;
        1486: data_ff <= 24'd300;
        1487: data_ff <= -24'd39;
        1488: data_ff <= 24'd6171221;
        1489: data_ff <= -24'd1735638;
        1490: data_ff <= 24'd931210;
        1491: data_ff <= -24'd575683;
        1492: data_ff <= 24'd371074;
        1493: data_ff <= -24'd239796;
        1494: data_ff <= 24'd152114;
        1495: data_ff <= -24'd93371;
        1496: data_ff <= 24'd54796;
        1497: data_ff <= -24'd30375;
        1498: data_ff <= 24'd15682;
        1499: data_ff <= -24'd7402;
        1500: data_ff <= 24'd3110;
        1501: data_ff <= -24'd1110;
        1502: data_ff <= 24'd301;
        1503: data_ff <= -24'd40;
        1504: data_ff <= 24'd6231246;
        1505: data_ff <= -24'd1734045;
        1506: data_ff <= 24'd928775;
        1507: data_ff <= -24'd573822;
        1508: data_ff <= 24'd369777;
        1509: data_ff <= -24'd238936;
        1510: data_ff <= 24'd151569;
        1511: data_ff <= -24'd93045;
        1512: data_ff <= 24'd54613;
        1513: data_ff <= -24'd30281;
        1514: data_ff <= 24'd15639;
        1515: data_ff <= -24'd7386;
        1516: data_ff <= 24'd3105;
        1517: data_ff <= -24'd1109;
        1518: data_ff <= 24'd301;
        1519: data_ff <= -24'd40;
        1520: data_ff <= 24'd6290684;
        1521: data_ff <= -24'd1731759;
        1522: data_ff <= 24'd925960;
        1523: data_ff <= -24'd571727;
        1524: data_ff <= 24'd368329;
        1525: data_ff <= -24'd237976;
        1526: data_ff <= 24'd150962;
        1527: data_ff <= -24'd92680;
        1528: data_ff <= 24'd54408;
        1529: data_ff <= -24'd30174;
        1530: data_ff <= 24'd15589;
        1531: data_ff <= -24'd7365;
        1532: data_ff <= 24'd3099;
        1533: data_ff <= -24'd1108;
        1534: data_ff <= 24'd302;
        1535: data_ff <= -24'd41;
        1536: data_ff <= 24'd6349522;
        1537: data_ff <= -24'd1728774;
        1538: data_ff <= 24'd922765;
        1539: data_ff <= -24'd569395;
        1540: data_ff <= 24'd366728;
        1541: data_ff <= -24'd236918;
        1542: data_ff <= 24'd150291;
        1543: data_ff <= -24'd92276;
        1544: data_ff <= 24'd54179;
        1545: data_ff <= -24'd30054;
        1546: data_ff <= 24'd15532;
        1547: data_ff <= -24'd7342;
        1548: data_ff <= 24'd3091;
        1549: data_ff <= -24'd1107;
        1550: data_ff <= 24'd302;
        1551: data_ff <= -24'd41;
        1552: data_ff <= 24'd6407746;
        1553: data_ff <= -24'd1725082;
        1554: data_ff <= 24'd919189;
        1555: data_ff <= -24'd566828;
        1556: data_ff <= 24'd364974;
        1557: data_ff <= -24'd235761;
        1558: data_ff <= 24'd149558;
        1559: data_ff <= -24'd91833;
        1560: data_ff <= 24'd53927;
        1561: data_ff <= -24'd29922;
        1562: data_ff <= 24'd15468;
        1563: data_ff <= -24'd7315;
        1564: data_ff <= 24'd3082;
        1565: data_ff <= -24'd1105;
        1566: data_ff <= 24'd302;
        1567: data_ff <= -24'd41;
        1568: data_ff <= 24'd6465344;
        1569: data_ff <= -24'd1720681;
        1570: data_ff <= 24'd915229;
        1571: data_ff <= -24'd564025;
        1572: data_ff <= 24'd363068;
        1573: data_ff <= -24'd234505;
        1574: data_ff <= 24'd148761;
        1575: data_ff <= -24'd91350;
        1576: data_ff <= 24'd53651;
        1577: data_ff <= -24'd29776;
        1578: data_ff <= 24'd15398;
        1579: data_ff <= -24'd7285;
        1580: data_ff <= 24'd3071;
        1581: data_ff <= -24'd1102;
        1582: data_ff <= 24'd302;
        1583: data_ff <= -24'd42;
        1584: data_ff <= 24'd6522301;
        1585: data_ff <= -24'd1715562;
        1586: data_ff <= 24'd910886;
        1587: data_ff <= -24'd560985;
        1588: data_ff <= 24'd361010;
        1589: data_ff <= -24'd233150;
        1590: data_ff <= 24'd147900;
        1591: data_ff <= -24'd90829;
        1592: data_ff <= 24'd53353;
        1593: data_ff <= -24'd29617;
        1594: data_ff <= 24'd15321;
        1595: data_ff <= -24'd7252;
        1596: data_ff <= 24'd3059;
        1597: data_ff <= -24'd1099;
        1598: data_ff <= 24'd302;
        1599: data_ff <= -24'd42;
        1600: data_ff <= 24'd6578605;
        1601: data_ff <= -24'd1709722;
        1602: data_ff <= 24'd906158;
        1603: data_ff <= -24'd557709;
        1604: data_ff <= 24'd358799;
        1605: data_ff <= -24'd231696;
        1606: data_ff <= 24'd146976;
        1607: data_ff <= -24'd90267;
        1608: data_ff <= 24'd53031;
        1609: data_ff <= -24'd29444;
        1610: data_ff <= 24'd15236;
        1611: data_ff <= -24'd7215;
        1612: data_ff <= 24'd3046;
        1613: data_ff <= -24'd1095;
        1614: data_ff <= 24'd302;
        1615: data_ff <= -24'd42;
        1616: data_ff <= 24'd6634243;
        1617: data_ff <= -24'd1703156;
        1618: data_ff <= 24'd901044;
        1619: data_ff <= -24'd554196;
        1620: data_ff <= 24'd356435;
        1621: data_ff <= -24'd230142;
        1622: data_ff <= 24'd145989;
        1623: data_ff <= -24'd89667;
        1624: data_ff <= 24'd52685;
        1625: data_ff <= -24'd29259;
        1626: data_ff <= 24'd15145;
        1627: data_ff <= -24'd7175;
        1628: data_ff <= 24'd3031;
        1629: data_ff <= -24'd1091;
        1630: data_ff <= 24'd301;
        1631: data_ff <= -24'd42;
        1632: data_ff <= 24'd6689202;
        1633: data_ff <= -24'd1695858;
        1634: data_ff <= 24'd895544;
        1635: data_ff <= -24'd550446;
        1636: data_ff <= 24'd353918;
        1637: data_ff <= -24'd228490;
        1638: data_ff <= 24'd144938;
        1639: data_ff <= -24'd89027;
        1640: data_ff <= 24'd52316;
        1641: data_ff <= -24'd29060;
        1642: data_ff <= 24'd15047;
        1643: data_ff <= -24'd7132;
        1644: data_ff <= 24'd3014;
        1645: data_ff <= -24'd1086;
        1646: data_ff <= 24'd300;
        1647: data_ff <= -24'd42;
        1648: data_ff <= 24'd6743469;
        1649: data_ff <= -24'd1687823;
        1650: data_ff <= 24'd889658;
        1651: data_ff <= -24'd546459;
        1652: data_ff <= 24'd351250;
        1653: data_ff <= -24'd226738;
        1654: data_ff <= 24'd143824;
        1655: data_ff <= -24'd88348;
        1656: data_ff <= 24'd51924;
        1657: data_ff <= -24'd28848;
        1658: data_ff <= 24'd14942;
        1659: data_ff <= -24'd7085;
        1660: data_ff <= 24'd2996;
        1661: data_ff <= -24'd1081;
        1662: data_ff <= 24'd299;
        1663: data_ff <= -24'd43;
        1664: data_ff <= 24'd6797032;
        1665: data_ff <= -24'd1679048;
        1666: data_ff <= 24'd883384;
        1667: data_ff <= -24'd542237;
        1668: data_ff <= 24'd348429;
        1669: data_ff <= -24'd224888;
        1670: data_ff <= 24'd142647;
        1671: data_ff <= -24'd87630;
        1672: data_ff <= 24'd51508;
        1673: data_ff <= -24'd28623;
        1674: data_ff <= 24'd14829;
        1675: data_ff <= -24'd7035;
        1676: data_ff <= 24'd2977;
        1677: data_ff <= -24'd1075;
        1678: data_ff <= 24'd298;
        1679: data_ff <= -24'd43;
        1680: data_ff <= 24'd6849878;
        1681: data_ff <= -24'd1669527;
        1682: data_ff <= 24'd876724;
        1683: data_ff <= -24'd537778;
        1684: data_ff <= 24'd345456;
        1685: data_ff <= -24'd222939;
        1686: data_ff <= 24'd141407;
        1687: data_ff <= -24'd86872;
        1688: data_ff <= 24'd51069;
        1689: data_ff <= -24'd28384;
        1690: data_ff <= 24'd14710;
        1691: data_ff <= -24'd6981;
        1692: data_ff <= 24'd2956;
        1693: data_ff <= -24'd1068;
        1694: data_ff <= 24'd297;
        1695: data_ff <= -24'd43;
        1696: data_ff <= 24'd6901996;
        1697: data_ff <= -24'd1659257;
        1698: data_ff <= 24'd869677;
        1699: data_ff <= -24'd533084;
        1700: data_ff <= 24'd342332;
        1701: data_ff <= -24'd220892;
        1702: data_ff <= 24'd140103;
        1703: data_ff <= -24'd86075;
        1704: data_ff <= 24'd50606;
        1705: data_ff <= -24'd28133;
        1706: data_ff <= 24'd14584;
        1707: data_ff <= -24'd6924;
        1708: data_ff <= 24'd2934;
        1709: data_ff <= -24'd1061;
        1710: data_ff <= 24'd296;
        1711: data_ff <= -24'd43;
        1712: data_ff <= 24'd6953372;
        1713: data_ff <= -24'd1648233;
        1714: data_ff <= 24'd862242;
        1715: data_ff <= -24'd528154;
        1716: data_ff <= 24'd339057;
        1717: data_ff <= -24'd218746;
        1718: data_ff <= 24'd138737;
        1719: data_ff <= -24'd85239;
        1720: data_ff <= 24'd50120;
        1721: data_ff <= -24'd27868;
        1722: data_ff <= 24'd14450;
        1723: data_ff <= -24'd6864;
        1724: data_ff <= 24'd2910;
        1725: data_ff <= -24'd1054;
        1726: data_ff <= 24'd294;
        1727: data_ff <= -24'd43;
        1728: data_ff <= 24'd7003996;
        1729: data_ff <= -24'd1636452;
        1730: data_ff <= 24'd854420;
        1731: data_ff <= -24'd522990;
        1732: data_ff <= 24'd335631;
        1733: data_ff <= -24'd216503;
        1734: data_ff <= 24'd137308;
        1735: data_ff <= -24'd84364;
        1736: data_ff <= 24'd49611;
        1737: data_ff <= -24'd27589;
        1738: data_ff <= 24'd14310;
        1739: data_ff <= -24'd6800;
        1740: data_ff <= 24'd2885;
        1741: data_ff <= -24'd1046;
        1742: data_ff <= 24'd293;
        1743: data_ff <= -24'd43;
        1744: data_ff <= 24'd7053856;
        1745: data_ff <= -24'd1623911;
        1746: data_ff <= 24'd846212;
        1747: data_ff <= -24'd517592;
        1748: data_ff <= 24'd332055;
        1749: data_ff <= -24'd214163;
        1750: data_ff <= 24'd135816;
        1751: data_ff <= -24'd83449;
        1752: data_ff <= 24'd49078;
        1753: data_ff <= -24'd27298;
        1754: data_ff <= 24'd14163;
        1755: data_ff <= -24'd6732;
        1756: data_ff <= 24'd2858;
        1757: data_ff <= -24'd1037;
        1758: data_ff <= 24'd291;
        1759: data_ff <= -24'd43;
        1760: data_ff <= 24'd7102939;
        1761: data_ff <= -24'd1610605;
        1762: data_ff <= 24'd837618;
        1763: data_ff <= -24'd511961;
        1764: data_ff <= 24'd328330;
        1765: data_ff <= -24'd211725;
        1766: data_ff <= 24'd134263;
        1767: data_ff <= -24'd82496;
        1768: data_ff <= 24'd48522;
        1769: data_ff <= -24'd26993;
        1770: data_ff <= 24'd14008;
        1771: data_ff <= -24'd6662;
        1772: data_ff <= 24'd2829;
        1773: data_ff <= -24'd1028;
        1774: data_ff <= 24'd289;
        1775: data_ff <= -24'd43;
        1776: data_ff <= 24'd7151235;
        1777: data_ff <= -24'd1596531;
        1778: data_ff <= 24'd828639;
        1779: data_ff <= -24'd506098;
        1780: data_ff <= 24'd324456;
        1781: data_ff <= -24'd209191;
        1782: data_ff <= 24'd132647;
        1783: data_ff <= -24'd81505;
        1784: data_ff <= 24'd47943;
        1785: data_ff <= -24'd26675;
        1786: data_ff <= 24'd13847;
        1787: data_ff <= -24'd6587;
        1788: data_ff <= 24'd2799;
        1789: data_ff <= -24'd1018;
        1790: data_ff <= 24'd287;
        1791: data_ff <= -24'd43;
        1792: data_ff <= 24'd7198732;
        1793: data_ff <= -24'd1581687;
        1794: data_ff <= 24'd819276;
        1795: data_ff <= -24'd500003;
        1796: data_ff <= 24'd320433;
        1797: data_ff <= -24'd206560;
        1798: data_ff <= 24'd130969;
        1799: data_ff <= -24'd80474;
        1800: data_ff <= 24'd47340;
        1801: data_ff <= -24'd26344;
        1802: data_ff <= 24'd13678;
        1803: data_ff <= -24'd6510;
        1804: data_ff <= 24'd2768;
        1805: data_ff <= -24'd1007;
        1806: data_ff <= 24'd284;
        1807: data_ff <= -24'd43;
        1808: data_ff <= 24'd7245419;
        1809: data_ff <= -24'd1566070;
        1810: data_ff <= 24'd809529;
        1811: data_ff <= -24'd493678;
        1812: data_ff <= 24'd316264;
        1813: data_ff <= -24'd203834;
        1814: data_ff <= 24'd129230;
        1815: data_ff <= -24'd79406;
        1816: data_ff <= 24'd46715;
        1817: data_ff <= -24'd25999;
        1818: data_ff <= 24'd13503;
        1819: data_ff <= -24'd6428;
        1820: data_ff <= 24'd2735;
        1821: data_ff <= -24'd996;
        1822: data_ff <= 24'd282;
        1823: data_ff <= -24'd43;
        1824: data_ff <= 24'd7291285;
        1825: data_ff <= -24'd1549676;
        1826: data_ff <= 24'd799399;
        1827: data_ff <= -24'd487124;
        1828: data_ff <= 24'd311948;
        1829: data_ff <= -24'd201013;
        1830: data_ff <= 24'd127430;
        1831: data_ff <= -24'd78299;
        1832: data_ff <= 24'd46066;
        1833: data_ff <= -24'd25642;
        1834: data_ff <= 24'd13320;
        1835: data_ff <= -24'd6344;
        1836: data_ff <= 24'd2700;
        1837: data_ff <= -24'd984;
        1838: data_ff <= 24'd279;
        1839: data_ff <= -24'd43;
        1840: data_ff <= 24'd7336320;
        1841: data_ff <= -24'd1532504;
        1842: data_ff <= 24'd788888;
        1843: data_ff <= -24'd480343;
        1844: data_ff <= 24'd307486;
        1845: data_ff <= -24'd198097;
        1846: data_ff <= 24'd125570;
        1847: data_ff <= -24'd77154;
        1848: data_ff <= 24'd45395;
        1849: data_ff <= -24'd25271;
        1850: data_ff <= 24'd13130;
        1851: data_ff <= -24'd6255;
        1852: data_ff <= 24'd2664;
        1853: data_ff <= -24'd972;
        1854: data_ff <= 24'd276;
        1855: data_ff <= -24'd43;
        1856: data_ff <= 24'd7380514;
        1857: data_ff <= -24'd1514551;
        1858: data_ff <= 24'd777998;
        1859: data_ff <= -24'd473334;
        1860: data_ff <= 24'd302879;
        1861: data_ff <= -24'd195088;
        1862: data_ff <= 24'd123649;
        1863: data_ff <= -24'd75971;
        1864: data_ff <= 24'd44701;
        1865: data_ff <= -24'd24888;
        1866: data_ff <= 24'd12934;
        1867: data_ff <= -24'd6164;
        1868: data_ff <= 24'd2626;
        1869: data_ff <= -24'd959;
        1870: data_ff <= 24'd273;
        1871: data_ff <= -24'd42;
        1872: data_ff <= 24'd7423855;
        1873: data_ff <= -24'd1495816;
        1874: data_ff <= 24'd766729;
        1875: data_ff <= -24'd466101;
        1876: data_ff <= 24'd298129;
        1877: data_ff <= -24'd191985;
        1878: data_ff <= 24'd121668;
        1879: data_ff <= -24'd74751;
        1880: data_ff <= 24'd43984;
        1881: data_ff <= -24'd24491;
        1882: data_ff <= 24'd12730;
        1883: data_ff <= -24'd6069;
        1884: data_ff <= 24'd2587;
        1885: data_ff <= -24'd946;
        1886: data_ff <= 24'd269;
        1887: data_ff <= -24'd42;
        1888: data_ff <= 24'd7466334;
        1889: data_ff <= -24'd1476296;
        1890: data_ff <= 24'd755084;
        1891: data_ff <= -24'd458644;
        1892: data_ff <= 24'd293237;
        1893: data_ff <= -24'd188790;
        1894: data_ff <= 24'd119627;
        1895: data_ff <= -24'd73494;
        1896: data_ff <= 24'd43245;
        1897: data_ff <= -24'd24082;
        1898: data_ff <= 24'd12520;
        1899: data_ff <= -24'd5970;
        1900: data_ff <= 24'd2546;
        1901: data_ff <= -24'd931;
        1902: data_ff <= 24'd266;
        1903: data_ff <= -24'd42;
        1904: data_ff <= 24'd7507940;
        1905: data_ff <= -24'd1455989;
        1906: data_ff <= 24'd743065;
        1907: data_ff <= -24'd450964;
        1908: data_ff <= 24'd288203;
        1909: data_ff <= -24'd185503;
        1910: data_ff <= 24'd117528;
        1911: data_ff <= -24'd72199;
        1912: data_ff <= 24'd42484;
        1913: data_ff <= -24'd23660;
        1914: data_ff <= 24'd12302;
        1915: data_ff <= -24'd5868;
        1916: data_ff <= 24'd2504;
        1917: data_ff <= -24'd917;
        1918: data_ff <= 24'd262;
        1919: data_ff <= -24'd41;
        1920: data_ff <= 24'd7548665;
        1921: data_ff <= -24'd1434895;
        1922: data_ff <= 24'd730672;
        1923: data_ff <= -24'd443065;
        1924: data_ff <= 24'd283028;
        1925: data_ff <= -24'd182125;
        1926: data_ff <= 24'd115370;
        1927: data_ff <= -24'd70868;
        1928: data_ff <= 24'd41700;
        1929: data_ff <= -24'd23225;
        1930: data_ff <= 24'd12078;
        1931: data_ff <= -24'd5763;
        1932: data_ff <= 24'd2460;
        1933: data_ff <= -24'd901;
        1934: data_ff <= 24'd258;
        1935: data_ff <= -24'd41;
        1936: data_ff <= 24'd7588498;
        1937: data_ff <= -24'd1413013;
        1938: data_ff <= 24'd717909;
        1939: data_ff <= -24'd434947;
        1940: data_ff <= 24'd277715;
        1941: data_ff <= -24'd178657;
        1942: data_ff <= 24'd113154;
        1943: data_ff <= -24'd69501;
        1944: data_ff <= 24'd40894;
        1945: data_ff <= -24'd22777;
        1946: data_ff <= 24'd11847;
        1947: data_ff <= -24'd5654;
        1948: data_ff <= 24'd2415;
        1949: data_ff <= -24'd886;
        1950: data_ff <= 24'd254;
        1951: data_ff <= -24'd41;
        1952: data_ff <= 24'd7627430;
        1953: data_ff <= -24'd1390340;
        1954: data_ff <= 24'd704778;
        1955: data_ff <= -24'd426613;
        1956: data_ff <= 24'd272265;
        1957: data_ff <= -24'd175099;
        1958: data_ff <= 24'd110880;
        1959: data_ff <= -24'd68097;
        1960: data_ff <= 24'd40067;
        1961: data_ff <= -24'd22317;
        1962: data_ff <= 24'd11609;
        1963: data_ff <= -24'd5542;
        1964: data_ff <= 24'd2368;
        1965: data_ff <= -24'd869;
        1966: data_ff <= 24'd250;
        1967: data_ff <= -24'd40;
        1968: data_ff <= 24'd7665452;
        1969: data_ff <= -24'd1366877;
        1970: data_ff <= 24'd691281;
        1971: data_ff <= -24'd418064;
        1972: data_ff <= 24'd266678;
        1973: data_ff <= -24'd171454;
        1974: data_ff <= 24'd108550;
        1975: data_ff <= -24'd66657;
        1976: data_ff <= 24'd39218;
        1977: data_ff <= -24'd21844;
        1978: data_ff <= 24'd11364;
        1979: data_ff <= -24'd5426;
        1980: data_ff <= 24'd2320;
        1981: data_ff <= -24'd852;
        1982: data_ff <= 24'd245;
        1983: data_ff <= -24'd40;
        1984: data_ff <= 24'd7702555;
        1985: data_ff <= -24'd1342623;
        1986: data_ff <= 24'd677421;
        1987: data_ff <= -24'd409303;
        1988: data_ff <= 24'd260956;
        1989: data_ff <= -24'd167721;
        1990: data_ff <= 24'd106164;
        1991: data_ff <= -24'd65183;
        1992: data_ff <= 24'd38347;
        1993: data_ff <= -24'd21359;
        1994: data_ff <= 24'd11112;
        1995: data_ff <= -24'd5307;
        1996: data_ff <= 24'd2270;
        1997: data_ff <= -24'd834;
        1998: data_ff <= 24'd240;
        1999: data_ff <= -24'd39;
        2000: data_ff <= 24'd7738730;
        2001: data_ff <= -24'd1317577;
        2002: data_ff <= 24'd663201;
        2003: data_ff <= -24'd400331;
        2004: data_ff <= 24'd255101;
        2005: data_ff <= -24'd163901;
        2006: data_ff <= 24'd103721;
        2007: data_ff <= -24'd63673;
        2008: data_ff <= 24'd37455;
        2009: data_ff <= -24'd20862;
        2010: data_ff <= 24'd10854;
        2011: data_ff <= -24'd5185;
        2012: data_ff <= 24'd2218;
        2013: data_ff <= -24'd816;
        2014: data_ff <= 24'd235;
        2015: data_ff <= -24'd38;
        2016: data_ff <= 24'd7773969;
        2017: data_ff <= -24'd1291739;
        2018: data_ff <= 24'd648623;
        2019: data_ff <= -24'd391151;
        2020: data_ff <= 24'd249114;
        2021: data_ff <= -24'd159997;
        2022: data_ff <= 24'd101224;
        2023: data_ff <= -24'd62128;
        2024: data_ff <= 24'd36542;
        2025: data_ff <= -24'd20352;
        2026: data_ff <= 24'd10590;
        2027: data_ff <= -24'd5059;
        2028: data_ff <= 24'd2165;
        2029: data_ff <= -24'd797;
        2030: data_ff <= 24'd230;
        2031: data_ff <= -24'd38;
        2032: data_ff <= 24'd7808264;
        2033: data_ff <= -24'd1265110;
        2034: data_ff <= 24'd633691;
        2035: data_ff <= -24'd381766;
        2036: data_ff <= 24'd242998;
        2037: data_ff <= -24'd156008;
        2038: data_ff <= 24'd98672;
        2039: data_ff <= -24'd60549;
        2040: data_ff <= 24'd35608;
        2041: data_ff <= -24'd19831;
        2042: data_ff <= 24'd10318;
        2043: data_ff <= -24'd4930;
        2044: data_ff <= 24'd2110;
        2045: data_ff <= -24'd777;
        2046: data_ff <= 24'd225;
        2047: data_ff <= -24'd37;
        2048: data_ff <= 24'd7841606;
        2049: data_ff <= -24'd1237690;
        2050: data_ff <= 24'd618407;
        2051: data_ff <= -24'd372177;
        2052: data_ff <= 24'd236753;
        2053: data_ff <= -24'd151936;
        2054: data_ff <= 24'd96067;
        2055: data_ff <= -24'd58937;
        2056: data_ff <= 24'd34654;
        2057: data_ff <= -24'd19297;
        2058: data_ff <= 24'd10040;
        2059: data_ff <= -24'd4798;
        2060: data_ff <= 24'd2054;
        2061: data_ff <= -24'd757;
        2062: data_ff <= 24'd219;
        2063: data_ff <= -24'd36;
        2064: data_ff <= 24'd7873988;
        2065: data_ff <= -24'd1209478;
        2066: data_ff <= 24'd602775;
        2067: data_ff <= -24'd362388;
        2068: data_ff <= 24'd230381;
        2069: data_ff <= -24'd147781;
        2070: data_ff <= 24'd93409;
        2071: data_ff <= -24'd57291;
        2072: data_ff <= 24'd33679;
        2073: data_ff <= -24'd18752;
        2074: data_ff <= 24'd9756;
        2075: data_ff <= -24'd4662;
        2076: data_ff <= 24'd1997;
        2077: data_ff <= -24'd736;
        2078: data_ff <= 24'd214;
        2079: data_ff <= -24'd36;
        2080: data_ff <= 24'd7905402;
        2081: data_ff <= -24'd1180477;
        2082: data_ff <= 24'd586799;
        2083: data_ff <= -24'd352401;
        2084: data_ff <= 24'd223885;
        2085: data_ff <= -24'd143547;
        2086: data_ff <= 24'd90699;
        2087: data_ff <= -24'd55612;
        2088: data_ff <= 24'd32684;
        2089: data_ff <= -24'd18195;
        2090: data_ff <= 24'd9465;
        2091: data_ff <= -24'd4523;
        2092: data_ff <= 24'd1937;
        2093: data_ff <= -24'd715;
        2094: data_ff <= 24'd208;
        2095: data_ff <= -24'd35;
        2096: data_ff <= 24'd7935840;
        2097: data_ff <= -24'd1150687;
        2098: data_ff <= 24'd570482;
        2099: data_ff <= -24'd342218;
        2100: data_ff <= 24'd217266;
        2101: data_ff <= -24'd139232;
        2102: data_ff <= 24'd87937;
        2103: data_ff <= -24'd53900;
        2104: data_ff <= 24'd31670;
        2105: data_ff <= -24'd17626;
        2106: data_ff <= 24'd9168;
        2107: data_ff <= -24'd4381;
        2108: data_ff <= 24'd1877;
        2109: data_ff <= -24'd693;
        2110: data_ff <= 24'd202;
        2111: data_ff <= -24'd34;
        2112: data_ff <= 24'd7965296;
        2113: data_ff <= -24'd1120108;
        2114: data_ff <= 24'd553829;
        2115: data_ff <= -24'd331843;
        2116: data_ff <= 24'd210525;
        2117: data_ff <= -24'd134839;
        2118: data_ff <= 24'd85124;
        2119: data_ff <= -24'd52157;
        2120: data_ff <= 24'd30636;
        2121: data_ff <= -24'd17046;
        2122: data_ff <= 24'd8865;
        2123: data_ff <= -24'd4236;
        2124: data_ff <= 24'd1815;
        2125: data_ff <= -24'd670;
        2126: data_ff <= 24'd195;
        2127: data_ff <= -24'd33;
        2128: data_ff <= 24'd7993762;
        2129: data_ff <= -24'd1088743;
        2130: data_ff <= 24'd536842;
        2131: data_ff <= -24'd321278;
        2132: data_ff <= 24'd203666;
        2133: data_ff <= -24'd130369;
        2134: data_ff <= 24'd82262;
        2135: data_ff <= -24'd50382;
        2136: data_ff <= 24'd29582;
        2137: data_ff <= -24'd16455;
        2138: data_ff <= 24'd8555;
        2139: data_ff <= -24'd4087;
        2140: data_ff <= 24'd1751;
        2141: data_ff <= -24'd647;
        2142: data_ff <= 24'd189;
        2143: data_ff <= -24'd32;
        2144: data_ff <= 24'd8021232;
        2145: data_ff <= -24'd1056594;
        2146: data_ff <= 24'd519526;
        2147: data_ff <= -24'd310527;
        2148: data_ff <= 24'd196690;
        2149: data_ff <= -24'd125823;
        2150: data_ff <= 24'd79351;
        2151: data_ff <= -24'd48576;
        2152: data_ff <= 24'd28510;
        2153: data_ff <= -24'd15853;
        2154: data_ff <= 24'd8240;
        2155: data_ff <= -24'd3936;
        2156: data_ff <= 24'd1686;
        2157: data_ff <= -24'd623;
        2158: data_ff <= 24'd182;
        2159: data_ff <= -24'd31;
        2160: data_ff <= 24'd8047699;
        2161: data_ff <= -24'd1023661;
        2162: data_ff <= 24'd501885;
        2163: data_ff <= -24'd299592;
        2164: data_ff <= 24'd189599;
        2165: data_ff <= -24'd121204;
        2166: data_ff <= 24'd76392;
        2167: data_ff <= -24'd46739;
        2168: data_ff <= 24'd27419;
        2169: data_ff <= -24'd15239;
        2170: data_ff <= 24'd7918;
        2171: data_ff <= -24'd3781;
        2172: data_ff <= 24'd1620;
        2173: data_ff <= -24'd598;
        2174: data_ff <= 24'd175;
        2175: data_ff <= -24'd30;
        2176: data_ff <= 24'd8073157;
        2177: data_ff <= -24'd989947;
        2178: data_ff <= 24'd483924;
        2179: data_ff <= -24'd288477;
        2180: data_ff <= 24'd182395;
        2181: data_ff <= -24'd116511;
        2182: data_ff <= 24'd73386;
        2183: data_ff <= -24'd44873;
        2184: data_ff <= 24'd26309;
        2185: data_ff <= -24'd14615;
        2186: data_ff <= 24'd7591;
        2187: data_ff <= -24'd3623;
        2188: data_ff <= 24'd1552;
        2189: data_ff <= -24'd573;
        2190: data_ff <= 24'd168;
        2191: data_ff <= -24'd29;
        2192: data_ff <= 24'd8097600;
        2193: data_ff <= -24'd955454;
        2194: data_ff <= 24'd465647;
        2195: data_ff <= -24'd277185;
        2196: data_ff <= 24'd175080;
        2197: data_ff <= -24'd111747;
        2198: data_ff <= 24'd70334;
        2199: data_ff <= -24'd42977;
        2200: data_ff <= 24'd25182;
        2201: data_ff <= -24'd13981;
        2202: data_ff <= 24'd7257;
        2203: data_ff <= -24'd3463;
        2204: data_ff <= 24'd1483;
        2205: data_ff <= -24'd548;
        2206: data_ff <= 24'd160;
        2207: data_ff <= -24'd28;
        2208: data_ff <= 24'd8121023;
        2209: data_ff <= -24'd920184;
        2210: data_ff <= 24'd447058;
        2211: data_ff <= -24'd265719;
        2212: data_ff <= 24'd167658;
        2213: data_ff <= -24'd106912;
        2214: data_ff <= 24'd67236;
        2215: data_ff <= -24'd41053;
        2216: data_ff <= 24'd24036;
        2217: data_ff <= -24'd13336;
        2218: data_ff <= 24'd6918;
        2219: data_ff <= -24'd3299;
        2220: data_ff <= 24'd1412;
        2221: data_ff <= -24'd521;
        2222: data_ff <= 24'd153;
        2223: data_ff <= -24'd26;
        2224: data_ff <= 24'd8143419;
        2225: data_ff <= -24'd884142;
        2226: data_ff <= 24'd428164;
        2227: data_ff <= -24'd254083;
        2228: data_ff <= 24'd160129;
        2229: data_ff <= -24'd102010;
        2230: data_ff <= 24'd64094;
        2231: data_ff <= -24'd39100;
        2232: data_ff <= 24'd22874;
        2233: data_ff <= -24'd12680;
        2234: data_ff <= 24'd6573;
        2235: data_ff <= -24'd3132;
        2236: data_ff <= 24'd1340;
        2237: data_ff <= -24'd495;
        2238: data_ff <= 24'd145;
        2239: data_ff <= -24'd25;
        2240: data_ff <= 24'd8164783;
        2241: data_ff <= -24'd847328;
        2242: data_ff <= 24'd408968;
        2243: data_ff <= -24'd242280;
        2244: data_ff <= 24'd152497;
        2245: data_ff <= -24'd97040;
        2246: data_ff <= 24'd60908;
        2247: data_ff <= -24'd37120;
        2248: data_ff <= 24'd21694;
        2249: data_ff <= -24'd12015;
        2250: data_ff <= 24'd6222;
        2251: data_ff <= -24'd2963;
        2252: data_ff <= 24'd1266;
        2253: data_ff <= -24'd467;
        2254: data_ff <= 24'd137;
        2255: data_ff <= -24'd24;
        2256: data_ff <= 24'd8185111;
        2257: data_ff <= -24'd809747;
        2258: data_ff <= 24'd389475;
        2259: data_ff <= -24'd230314;
        2260: data_ff <= 24'd144763;
        2261: data_ff <= -24'd92005;
        2262: data_ff <= 24'd57681;
        2263: data_ff <= -24'd35113;
        2264: data_ff <= 24'd20498;
        2265: data_ff <= -24'd11340;
        2266: data_ff <= 24'd5866;
        2267: data_ff <= -24'd2790;
        2268: data_ff <= 24'd1191;
        2269: data_ff <= -24'd439;
        2270: data_ff <= 24'd129;
        2271: data_ff <= -24'd22;
        2272: data_ff <= 24'd8204397;
        2273: data_ff <= -24'd771402;
        2274: data_ff <= 24'd369692;
        2275: data_ff <= -24'd218188;
        2276: data_ff <= 24'd136931;
        2277: data_ff <= -24'd86907;
        2278: data_ff <= 24'd54412;
        2279: data_ff <= -24'd33079;
        2280: data_ff <= 24'd19286;
        2281: data_ff <= -24'd10655;
        2282: data_ff <= 24'd5505;
        2283: data_ff <= -24'd2615;
        2284: data_ff <= 24'd1115;
        2285: data_ff <= -24'd411;
        2286: data_ff <= 24'd120;
        2287: data_ff <= -24'd21;
        2288: data_ff <= 24'd8222636;
        2289: data_ff <= -24'd732296;
        2290: data_ff <= 24'd349623;
        2291: data_ff <= -24'd205907;
        2292: data_ff <= 24'd129003;
        2293: data_ff <= -24'd81747;
        2294: data_ff <= 24'd51103;
        2295: data_ff <= -24'd31020;
        2296: data_ff <= 24'd18057;
        2297: data_ff <= -24'd9961;
        2298: data_ff <= 24'd5138;
        2299: data_ff <= -24'd2437;
        2300: data_ff <= 24'd1038;
        2301: data_ff <= -24'd382;
        2302: data_ff <= 24'd112;
        2303: data_ff <= -24'd20;
        2304: data_ff <= 24'd8239826;
        2305: data_ff <= -24'd692433;
        2306: data_ff <= 24'd329273;
        2307: data_ff <= -24'd193473;
        2308: data_ff <= 24'd120982;
        2309: data_ff <= -24'd76526;
        2310: data_ff <= 24'd47754;
        2311: data_ff <= -24'd28936;
        2312: data_ff <= 24'd16813;
        2313: data_ff <= -24'd9257;
        2314: data_ff <= 24'd4766;
        2315: data_ff <= -24'd2256;
        2316: data_ff <= 24'd959;
        2317: data_ff <= -24'd352;
        2318: data_ff <= 24'd103;
        2319: data_ff <= -24'd18;
        2320: data_ff <= 24'd8255961;
        2321: data_ff <= -24'd651818;
        2322: data_ff <= 24'd308649;
        2323: data_ff <= -24'd180892;
        2324: data_ff <= 24'd112869;
        2325: data_ff <= -24'd71247;
        2326: data_ff <= 24'd44368;
        2327: data_ff <= -24'd26828;
        2328: data_ff <= 24'd15554;
        2329: data_ff <= -24'd8545;
        2330: data_ff <= 24'd4389;
        2331: data_ff <= -24'd2073;
        2332: data_ff <= 24'd879;
        2333: data_ff <= -24'd322;
        2334: data_ff <= 24'd94;
        2335: data_ff <= -24'd16;
        2336: data_ff <= 24'd8271038;
        2337: data_ff <= -24'd610454;
        2338: data_ff <= 24'd287756;
        2339: data_ff <= -24'd168167;
        2340: data_ff <= 24'd104668;
        2341: data_ff <= -24'd65910;
        2342: data_ff <= 24'd40945;
        2343: data_ff <= -24'd24695;
        2344: data_ff <= 24'd14281;
        2345: data_ff <= -24'd7824;
        2346: data_ff <= 24'd4007;
        2347: data_ff <= -24'd1887;
        2348: data_ff <= 24'd797;
        2349: data_ff <= -24'd291;
        2350: data_ff <= 24'd85;
        2351: data_ff <= -24'd15;
        2352: data_ff <= 24'd8285052;
        2353: data_ff <= -24'd568347;
        2354: data_ff <= 24'd266601;
        2355: data_ff <= -24'd155302;
        2356: data_ff <= 24'd96381;
        2357: data_ff <= -24'd60519;
        2358: data_ff <= 24'd37486;
        2359: data_ff <= -24'd22540;
        2360: data_ff <= 24'd12993;
        2361: data_ff <= -24'd7094;
        2362: data_ff <= 24'd3620;
        2363: data_ff <= -24'd1698;
        2364: data_ff <= 24'd715;
        2365: data_ff <= -24'd260;
        2366: data_ff <= 24'd75;
        2367: data_ff <= -24'd13;
        2368: data_ff <= 24'd8298002;
        2369: data_ff <= -24'd525500;
        2370: data_ff <= 24'd245189;
        2371: data_ff <= -24'd142301;
        2372: data_ff <= 24'd88012;
        2373: data_ff <= -24'd55075;
        2374: data_ff <= 24'd33993;
        2375: data_ff <= -24'd20363;
        2376: data_ff <= 24'd11691;
        2377: data_ff <= -24'd6356;
        2378: data_ff <= 24'd3229;
        2379: data_ff <= -24'd1507;
        2380: data_ff <= 24'd631;
        2381: data_ff <= -24'd228;
        2382: data_ff <= 24'd66;
        2383: data_ff <= -24'd11;
        2384: data_ff <= 24'd8309883;
        2385: data_ff <= -24'd481919;
        2386: data_ff <= 24'd223526;
        2387: data_ff <= -24'd129169;
        2388: data_ff <= 24'd79563;
        2389: data_ff <= -24'd49579;
        2390: data_ff <= 24'd30466;
        2391: data_ff <= -24'd18164;
        2392: data_ff <= 24'd10375;
        2393: data_ff <= -24'd5610;
        2394: data_ff <= 24'd2833;
        2395: data_ff <= -24'd1313;
        2396: data_ff <= 24'd546;
        2397: data_ff <= -24'd196;
        2398: data_ff <= 24'd56;
        2399: data_ff <= -24'd9;
        2400: data_ff <= 24'd8320693;
        2401: data_ff <= -24'd437608;
        2402: data_ff <= 24'd201619;
        2403: data_ff <= -24'd115910;
        2404: data_ff <= 24'd71037;
        2405: data_ff <= -24'd44034;
        2406: data_ff <= 24'd26907;
        2407: data_ff <= -24'd15945;
        2408: data_ff <= 24'd9047;
        2409: data_ff <= -24'd4856;
        2410: data_ff <= 24'd2432;
        2411: data_ff <= -24'd1117;
        2412: data_ff <= 24'd460;
        2413: data_ff <= -24'd163;
        2414: data_ff <= 24'd46;
        2415: data_ff <= -24'd8;
        2416: data_ff <= 24'd8330430;
        2417: data_ff <= -24'd392574;
        2418: data_ff <= 24'd179474;
        2419: data_ff <= -24'd102528;
        2420: data_ff <= 24'd62436;
        2421: data_ff <= -24'd38442;
        2422: data_ff <= 24'd23316;
        2423: data_ff <= -24'd13705;
        2424: data_ff <= 24'd7706;
        2425: data_ff <= -24'd4094;
        2426: data_ff <= 24'd2027;
        2427: data_ff <= -24'd919;
        2428: data_ff <= 24'd372;
        2429: data_ff <= -24'd130;
        2430: data_ff <= 24'd36;
        2431: data_ff <= -24'd6;
        2432: data_ff <= 24'd8339090;
        2433: data_ff <= -24'd346821;
        2434: data_ff <= 24'd157098;
        2435: data_ff <= -24'd89027;
        2436: data_ff <= 24'd53765;
        2437: data_ff <= -24'd32803;
        2438: data_ff <= 24'd19697;
        2439: data_ff <= -24'd11446;
        2440: data_ff <= 24'd6353;
        2441: data_ff <= -24'd3325;
        2442: data_ff <= 24'd1618;
        2443: data_ff <= -24'd719;
        2444: data_ff <= 24'd284;
        2445: data_ff <= -24'd96;
        2446: data_ff <= 24'd25;
        2447: data_ff <= -24'd4;
        2448: data_ff <= 24'd8346673;
        2449: data_ff <= -24'd300356;
        2450: data_ff <= 24'd134498;
        2451: data_ff <= -24'd75413;
        2452: data_ff <= 24'd45025;
        2453: data_ff <= -24'd27121;
        2454: data_ff <= 24'd16048;
        2455: data_ff <= -24'd9169;
        2456: data_ff <= 24'd4989;
        2457: data_ff <= -24'd2549;
        2458: data_ff <= 24'd1204;
        2459: data_ff <= -24'd516;
        2460: data_ff <= 24'd194;
        2461: data_ff <= -24'd62;
        2462: data_ff <= 24'd15;
        2463: data_ff <= -24'd2;
        2464: data_ff <= 24'd8353175;
        2465: data_ff <= -24'd253184;
        2466: data_ff <= 24'd111680;
        2467: data_ff <= -24'd61690;
        2468: data_ff <= 24'd36220;
        2469: data_ff <= -24'd21398;
        2470: data_ff <= 24'd12373;
        2471: data_ff <= -24'd6875;
        2472: data_ff <= 24'd3613;
        2473: data_ff <= -24'd1766;
        2474: data_ff <= 24'd787;
        2475: data_ff <= -24'd311;
        2476: data_ff <= 24'd104;
        2477: data_ff <= -24'd27;
        2478: data_ff <= 24'd4;
        2479: data_ff <= -24'd0;
        2480: data_ff <= 24'd8358596;
        2481: data_ff <= -24'd205312;
        2482: data_ff <= 24'd88651;
        2483: data_ff <= -24'd47862;
        2484: data_ff <= 24'd27353;
        2485: data_ff <= -24'd15635;
        2486: data_ff <= 24'd8672;
        2487: data_ff <= -24'd4563;
        2488: data_ff <= 24'd2226;
        2489: data_ff <= -24'd977;
        2490: data_ff <= 24'd366;
        2491: data_ff <= -24'd104;
        2492: data_ff <= 24'd12;
        2493: data_ff <= 24'd8;
        2494: data_ff <= -24'd6;
        2495: data_ff <= 24'd2;
        2496: data_ff <= 24'd8362935;
        2497: data_ff <= -24'd156746;
        2498: data_ff <= 24'd65419;
        2499: data_ff <= -24'd33934;
        2500: data_ff <= 24'd18427;
        2501: data_ff <= -24'd9834;
        2502: data_ff <= 24'd4946;
        2503: data_ff <= -24'd2235;
        2504: data_ff <= 24'd829;
        2505: data_ff <= -24'd181;
        2506: data_ff <= -24'd58;
        2507: data_ff <= 24'd104;
        2508: data_ff <= -24'd80;
        2509: data_ff <= 24'd43;
        2510: data_ff <= -24'd17;
        2511: data_ff <= 24'd4;
        2512: data_ff <= 24'd8366190;
        2513: data_ff <= -24'd107493;
        2514: data_ff <= 24'd41991;
        2515: data_ff <= -24'd19911;
        2516: data_ff <= 24'd9446;
        2517: data_ff <= -24'd3998;
        2518: data_ff <= 24'd1197;
        2519: data_ff <= 24'd106;
        2520: data_ff <= -24'd576;
        2521: data_ff <= 24'd619;
        2522: data_ff <= -24'd486;
        2523: data_ff <= 24'd315;
        2524: data_ff <= -24'd173;
        2525: data_ff <= 24'd79;
        2526: data_ff <= -24'd28;
        2527: data_ff <= 24'd6;
        2528: data_ff <= 24'd8368360;
        2529: data_ff <= -24'd57559;
        2530: data_ff <= 24'd18374;
        2531: data_ff <= -24'd5798;
        2532: data_ff <= 24'd411;
        2533: data_ff <= 24'd1871;
        2534: data_ff <= -24'd2573;
        2535: data_ff <= 24'd2463;
        2536: data_ff <= -24'd1992;
        2537: data_ff <= 24'd1427;
        2538: data_ff <= -24'd918;
        2539: data_ff <= 24'd528;
        2540: data_ff <= -24'd268;
        2541: data_ff <= 24'd116;
        2542: data_ff <= -24'd40;
        2543: data_ff <= 24'd8;
        2544: data_ff <= 24'd8369445;
        2545: data_ff <= -24'd6952;
        2546: data_ff <= -24'd5424;
        2547: data_ff <= 24'd8399;
        2548: data_ff <= -24'd8671;
        2549: data_ff <= 24'd7771;
        2550: data_ff <= -24'd6364;
        2551: data_ff <= 24'd4834;
        2552: data_ff <= -24'd3416;
        2553: data_ff <= 24'd2240;
        2554: data_ff <= -24'd1352;
        2555: data_ff <= 24'd743;
        2556: data_ff <= -24'd364;
        2557: data_ff <= 24'd153;
        2558: data_ff <= -24'd52;
        2559: data_ff <= 24'd11;

        default: data_ff <= 0;
    endcase
end
endmodule
