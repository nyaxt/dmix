// Polyphase filter bank for upsampling from 44100.0kHz to 48000.0kHz
// Depth: 32

module rom_firbank_441_480(
    input clk,
    input [11:0] addr,
    output [23:0] data);
reg [23:0] data_ff;
assign data = data_ff;
always @(posedge clk) begin
    case(addr)
        0: data_ff <= 24'h005690; // 22160
        1: data_ff <= 24'hFFC696; // -14698
        2: data_ff <= 24'h002C4B; // 11339
        3: data_ff <= 24'hFFDD3C; // -8900
        4: data_ff <= 24'h001AC2; // 6850
        5: data_ff <= 24'hFFEC21; // -5087
        6: data_ff <= 24'h000E18; // 3608
        7: data_ff <= 24'hFFF688; // -2424
        8: data_ff <= 24'h0005F9; // 1529
        9: data_ff <= 24'hFFFC81; // -895
        10: data_ff <= 24'h0001DF; // 479
        11: data_ff <= 24'hFFFF1A; // -230
        12: data_ff <= 24'h00005F; // 95
        13: data_ff <= 24'hFFFFE1; // -31
        14: data_ff <= 24'h000006; // 6
        15: data_ff <= 24'h000000; // 0
        16: data_ff <= 24'h00BBFD; // 48125
        17: data_ff <= 24'hFF9771; // -26767
        18: data_ff <= 24'h004854; // 18516
        19: data_ff <= 24'hFFCB52; // -13486
        20: data_ff <= 24'h002665; // 9829
        21: data_ff <= 24'hFFE4A7; // -7001
        22: data_ff <= 24'h0012C6; // 4806
        23: data_ff <= 24'hFFF3B8; // -3144
        24: data_ff <= 24'h000794; // 1940
        25: data_ff <= 24'hFFFBA5; // -1115
        26: data_ff <= 24'h00024C; // 588
        27: data_ff <= 24'hFFFEEA; // -278
        28: data_ff <= 24'h000072; // 114
        29: data_ff <= 24'hFFFFDB; // -37
        30: data_ff <= 24'h000008; // 8
        31: data_ff <= 24'h000000; // 0
        32: data_ff <= 24'h0122B1; // 74417
        33: data_ff <= 24'hFF67FC; // -38916
        34: data_ff <= 24'h006480; // 25728
        35: data_ff <= 24'hFFB954; // -18092
        36: data_ff <= 24'h003213; // 12819
        37: data_ff <= 24'hFFDD25; // -8923
        38: data_ff <= 24'h001779; // 6009
        39: data_ff <= 24'hFFF0E4; // -3868
        40: data_ff <= 24'h000932; // 2354
        41: data_ff <= 24'hFFFAC7; // -1337
        42: data_ff <= 24'h0002BA; // 698
        43: data_ff <= 24'hFFFEB8; // -328
        44: data_ff <= 24'h000085; // 133
        45: data_ff <= 24'hFFFFD5; // -43
        46: data_ff <= 24'h000009; // 9
        47: data_ff <= 24'h000000; // 0
        48: data_ff <= 24'h018AA5; // 101029
        49: data_ff <= 24'hFF383D; // -51139
        50: data_ff <= 24'h0080CC; // 32972
        51: data_ff <= 24'hFFA744; // -22716
        52: data_ff <= 24'h003DCD; // 15821
        53: data_ff <= 24'hFFD59B; // -10853
        54: data_ff <= 24'h001C30; // 7216
        55: data_ff <= 24'hFFEE0D; // -4595
        56: data_ff <= 24'h000AD2; // 2770
        57: data_ff <= 24'hFFF9E8; // -1560
        58: data_ff <= 24'h000329; // 809
        59: data_ff <= 24'hFFFE87; // -377
        60: data_ff <= 24'h000098; // 152
        61: data_ff <= 24'hFFFFCE; // -50
        62: data_ff <= 24'h00000A; // 10
        63: data_ff <= 24'h000000; // 0
        64: data_ff <= 24'h01F3D8; // 127960
        65: data_ff <= 24'hFF0836; // -63434
        66: data_ff <= 24'h009D37; // 40247
        67: data_ff <= 24'hFF9524; // -27356
        68: data_ff <= 24'h004991; // 18833
        69: data_ff <= 24'hFFCE0B; // -12789
        70: data_ff <= 24'h0020ED; // 8429
        71: data_ff <= 24'hFFEB33; // -5325
        72: data_ff <= 24'h000C73; // 3187
        73: data_ff <= 24'hFFF907; // -1785
        74: data_ff <= 24'h000398; // 920
        75: data_ff <= 24'hFFFE55; // -427
        76: data_ff <= 24'h0000AC; // 172
        77: data_ff <= 24'hFFFFC8; // -56
        78: data_ff <= 24'h00000B; // 11
        79: data_ff <= 24'hFFFFFF; // -1
        80: data_ff <= 24'h025E43; // 155203
        81: data_ff <= 24'hFED7EC; // -75796
        82: data_ff <= 24'h00B9BC; // 47548
        83: data_ff <= 24'hFF82F5; // -32011
        84: data_ff <= 24'h00555F; // 21855
        85: data_ff <= 24'hFFC674; // -14732
        86: data_ff <= 24'h0025AD; // 9645
        87: data_ff <= 24'hFFE856; // -6058
        88: data_ff <= 24'h000E17; // 3607
        89: data_ff <= 24'hFFF826; // -2010
        90: data_ff <= 24'h000408; // 1032
        91: data_ff <= 24'hFFFE23; // -477
        92: data_ff <= 24'h0000C0; // 192
        93: data_ff <= 24'hFFFFC2; // -62
        94: data_ff <= 24'h00000D; // 13
        95: data_ff <= 24'hFFFFFF; // -1
        96: data_ff <= 24'h02C9E4; // 182756
        97: data_ff <= 24'hFEA763; // -88221
        98: data_ff <= 24'h00D65A; // 54874
        99: data_ff <= 24'hFF70BA; // -36678
        100: data_ff <= 24'h006134; // 24884
        101: data_ff <= 24'hFFBED9; // -16679
        102: data_ff <= 24'h002A71; // 10865
        103: data_ff <= 24'hFFE577; // -6793
        104: data_ff <= 24'h000FBC; // 4028
        105: data_ff <= 24'hFFF743; // -2237
        106: data_ff <= 24'h000479; // 1145
        107: data_ff <= 24'hFFFDF0; // -528
        108: data_ff <= 24'h0000D4; // 212
        109: data_ff <= 24'hFFFFBB; // -69
        110: data_ff <= 24'h00000E; // 14
        111: data_ff <= 24'hFFFFFF; // -1
        112: data_ff <= 24'h0336B5; // 210613
        113: data_ff <= 24'hFE769F; // -100705
        114: data_ff <= 24'h00F30F; // 62223
        115: data_ff <= 24'hFF5E73; // -41357
        116: data_ff <= 24'h006D0F; // 27919
        117: data_ff <= 24'hFFB739; // -18631
        118: data_ff <= 24'h002F39; // 12089
        119: data_ff <= 24'hFFE296; // -7530
        120: data_ff <= 24'h001163; // 4451
        121: data_ff <= 24'hFFF660; // -2464
        122: data_ff <= 24'h0004EA; // 1258
        123: data_ff <= 24'hFFFDBD; // -579
        124: data_ff <= 24'h0000E8; // 232
        125: data_ff <= 24'hFFFFB5; // -75
        126: data_ff <= 24'h000010; // 16
        127: data_ff <= 24'hFFFFFF; // -1
        128: data_ff <= 24'h03A4B3; // 238771
        129: data_ff <= 24'hFE45A4; // -113244
        130: data_ff <= 24'h010FD6; // 69590
        131: data_ff <= 24'hFF4C23; // -46045
        132: data_ff <= 24'h0078F0; // 30960
        133: data_ff <= 24'hFFAF95; // -20587
        134: data_ff <= 24'h003403; // 13315
        135: data_ff <= 24'hFFDFB2; // -8270
        136: data_ff <= 24'h00130B; // 4875
        137: data_ff <= 24'hFFF57B; // -2693
        138: data_ff <= 24'h00055B; // 1371
        139: data_ff <= 24'hFFFD8A; // -630
        140: data_ff <= 24'h0000FC; // 252
        141: data_ff <= 24'hFFFFAE; // -82
        142: data_ff <= 24'h000011; // 17
        143: data_ff <= 24'hFFFFFF; // -1
        144: data_ff <= 24'h0413D8; // 267224
        145: data_ff <= 24'hFE1478; // -125832
        146: data_ff <= 24'h012CAE; // 76974
        147: data_ff <= 24'hFF39CC; // -50740
        148: data_ff <= 24'h0084D6; // 34006
        149: data_ff <= 24'hFFA7EE; // -22546
        150: data_ff <= 24'h0038CF; // 14543
        151: data_ff <= 24'hFFDCCD; // -9011
        152: data_ff <= 24'h0014B4; // 5300
        153: data_ff <= 24'hFFF496; // -2922
        154: data_ff <= 24'h0005CE; // 1486
        155: data_ff <= 24'hFFFD57; // -681
        156: data_ff <= 24'h000110; // 272
        157: data_ff <= 24'hFFFFA8; // -88
        158: data_ff <= 24'h000012; // 18
        159: data_ff <= 24'hFFFFFF; // -1
        160: data_ff <= 24'h048421; // 295969
        161: data_ff <= 24'hFDE31D; // -138467
        162: data_ff <= 24'h014994; // 84372
        163: data_ff <= 24'hFF276F; // -55441
        164: data_ff <= 24'h0090BF; // 37055
        165: data_ff <= 24'hFFA045; // -24507
        166: data_ff <= 24'h003D9C; // 15772
        167: data_ff <= 24'hFFD9E7; // -9753
        168: data_ff <= 24'h00165F; // 5727
        169: data_ff <= 24'hFFF3B0; // -3152
        170: data_ff <= 24'h000640; // 1600
        171: data_ff <= 24'hFFFD23; // -733
        172: data_ff <= 24'h000125; // 293
        173: data_ff <= 24'hFFFFA1; // -95
        174: data_ff <= 24'h000014; // 20
        175: data_ff <= 24'hFFFFFF; // -1
        176: data_ff <= 24'h04F588; // 325000
        177: data_ff <= 24'hFDB198; // -151144
        178: data_ff <= 24'h016684; // 91780
        179: data_ff <= 24'hFF150D; // -60147
        180: data_ff <= 24'h009CAA; // 40106
        181: data_ff <= 24'hFF989A; // -26470
        182: data_ff <= 24'h00426C; // 17004
        183: data_ff <= 24'hFFD700; // -10496
        184: data_ff <= 24'h00180A; // 6154
        185: data_ff <= 24'hFFF2CA; // -3382
        186: data_ff <= 24'h0006B3; // 1715
        187: data_ff <= 24'hFFFCEF; // -785
        188: data_ff <= 24'h000139; // 313
        189: data_ff <= 24'hFFFF9B; // -101
        190: data_ff <= 24'h000015; // 21
        191: data_ff <= 24'hFFFFFF; // -1
        192: data_ff <= 24'h056808; // 354312
        193: data_ff <= 24'hFD7FEF; // -163857
        194: data_ff <= 24'h01837D; // 99197
        195: data_ff <= 24'hFF02AA; // -64854
        196: data_ff <= 24'h00A895; // 43157
        197: data_ff <= 24'hFF90EF; // -28433
        198: data_ff <= 24'h00473B; // 18235
        199: data_ff <= 24'hFFD417; // -11241
        200: data_ff <= 24'h0019B6; // 6582
        201: data_ff <= 24'hFFF1E2; // -3614
        202: data_ff <= 24'h000727; // 1831
        203: data_ff <= 24'hFFFCBA; // -838
        204: data_ff <= 24'h00014E; // 334
        205: data_ff <= 24'hFFFF94; // -108
        206: data_ff <= 24'h000017; // 23
        207: data_ff <= 24'hFFFFFF; // -1
        208: data_ff <= 24'h05DB9D; // 383901
        209: data_ff <= 24'hFD4E24; // -176604
        210: data_ff <= 24'h01A07B; // 106619
        211: data_ff <= 24'hFEF047; // -69561
        212: data_ff <= 24'h00B481; // 46209
        213: data_ff <= 24'hFF8944; // -30396
        214: data_ff <= 24'h004C0C; // 19468
        215: data_ff <= 24'hFFD12F; // -11985
        216: data_ff <= 24'h001B62; // 7010
        217: data_ff <= 24'hFFF0FB; // -3845
        218: data_ff <= 24'h00079B; // 1947
        219: data_ff <= 24'hFFFC86; // -890
        220: data_ff <= 24'h000163; // 355
        221: data_ff <= 24'hFFFF8D; // -115
        222: data_ff <= 24'h000018; // 24
        223: data_ff <= 24'hFFFFFF; // -1
        224: data_ff <= 24'h065042; // 413762
        225: data_ff <= 24'hFD1C3E; // -189378
        226: data_ff <= 24'h01BD7C; // 114044
        227: data_ff <= 24'hFEDDE5; // -74267
        228: data_ff <= 24'h00C06A; // 49258
        229: data_ff <= 24'hFF819A; // -32358
        230: data_ff <= 24'h0050DB; // 20699
        231: data_ff <= 24'hFFCE46; // -12730
        232: data_ff <= 24'h001D0F; // 7439
        233: data_ff <= 24'hFFF013; // -4077
        234: data_ff <= 24'h00080F; // 2063
        235: data_ff <= 24'hFFFC51; // -943
        236: data_ff <= 24'h000178; // 376
        237: data_ff <= 24'hFFFF86; // -122
        238: data_ff <= 24'h00001A; // 26
        239: data_ff <= 24'hFFFFFE; // -2
        240: data_ff <= 24'h06C5F2; // 443890
        241: data_ff <= 24'hFCEA3F; // -202177
        242: data_ff <= 24'h01DA7C; // 121468
        243: data_ff <= 24'hFECB86; // -78970
        244: data_ff <= 24'h00CC51; // 52305
        245: data_ff <= 24'hFF79F1; // -34319
        246: data_ff <= 24'h0055AB; // 21931
        247: data_ff <= 24'hFFCB5D; // -13475
        248: data_ff <= 24'h001EBB; // 7867
        249: data_ff <= 24'hFFEF2B; // -4309
        250: data_ff <= 24'h000883; // 2179
        251: data_ff <= 24'hFFFC1C; // -996
        252: data_ff <= 24'h00018D; // 397
        253: data_ff <= 24'hFFFF7F; // -129
        254: data_ff <= 24'h00001C; // 28
        255: data_ff <= 24'hFFFFFE; // -2
        256: data_ff <= 24'h073CA6; // 474278
        257: data_ff <= 24'hFCB82E; // -214994
        258: data_ff <= 24'h01F77A; // 128890
        259: data_ff <= 24'hFEB92D; // -83667
        260: data_ff <= 24'h00D834; // 55348
        261: data_ff <= 24'hFF724B; // -36277
        262: data_ff <= 24'h005A79; // 23161
        263: data_ff <= 24'hFFC875; // -14219
        264: data_ff <= 24'h002068; // 8296
        265: data_ff <= 24'hFFEE43; // -4541
        266: data_ff <= 24'h0008F8; // 2296
        267: data_ff <= 24'hFFFBE7; // -1049
        268: data_ff <= 24'h0001A2; // 418
        269: data_ff <= 24'hFFFF78; // -136
        270: data_ff <= 24'h00001D; // 29
        271: data_ff <= 24'hFFFFFE; // -2
        272: data_ff <= 24'h07B45B; // 504923
        273: data_ff <= 24'hFC860E; // -227826
        274: data_ff <= 24'h021471; // 136305
        275: data_ff <= 24'hFEA6DB; // -88357
        276: data_ff <= 24'h00E412; // 58386
        277: data_ff <= 24'hFF6AA7; // -38233
        278: data_ff <= 24'h005F45; // 24389
        279: data_ff <= 24'hFFC58D; // -14963
        280: data_ff <= 24'h002215; // 8725
        281: data_ff <= 24'hFFED5A; // -4774
        282: data_ff <= 24'h00096C; // 2412
        283: data_ff <= 24'hFFFBB2; // -1102
        284: data_ff <= 24'h0001B7; // 439
        285: data_ff <= 24'hFFFF71; // -143
        286: data_ff <= 24'h00001F; // 31
        287: data_ff <= 24'hFFFFFE; // -2
        288: data_ff <= 24'h082D0B; // 535819
        289: data_ff <= 24'hFC53E4; // -240668
        290: data_ff <= 24'h02315F; // 143711
        291: data_ff <= 24'hFE9491; // -93039
        292: data_ff <= 24'h00EFEA; // 61418
        293: data_ff <= 24'hFF6308; // -40184
        294: data_ff <= 24'h00640F; // 25615
        295: data_ff <= 24'hFFC2A7; // -15705
        296: data_ff <= 24'h0023C1; // 9153
        297: data_ff <= 24'hFFEC72; // -5006
        298: data_ff <= 24'h0009E1; // 2529
        299: data_ff <= 24'hFFFB7D; // -1155
        300: data_ff <= 24'h0001CD; // 461
        301: data_ff <= 24'hFFFF6A; // -150
        302: data_ff <= 24'h000021; // 33
        303: data_ff <= 24'hFFFFFE; // -2
        304: data_ff <= 24'h08A6B0; // 566960
        305: data_ff <= 24'hFC21B5; // -253515
        306: data_ff <= 24'h024E41; // 151105
        307: data_ff <= 24'hFE8253; // -97709
        308: data_ff <= 24'h00FBB9; // 64441
        309: data_ff <= 24'hFF5B6E; // -42130
        310: data_ff <= 24'h0068D7; // 26839
        311: data_ff <= 24'hFFBFC1; // -16447
        312: data_ff <= 24'h00256D; // 9581
        313: data_ff <= 24'hFFEB8A; // -5238
        314: data_ff <= 24'h000A56; // 2646
        315: data_ff <= 24'hFFFB48; // -1208
        316: data_ff <= 24'h0001E2; // 482
        317: data_ff <= 24'hFFFF63; // -157
        318: data_ff <= 24'h000022; // 34
        319: data_ff <= 24'hFFFFFE; // -2
        320: data_ff <= 24'h092144; // 598340
        321: data_ff <= 24'hFBEF86; // -266362
        322: data_ff <= 24'h026B15; // 158485
        323: data_ff <= 24'hFE7021; // -102367
        324: data_ff <= 24'h010780; // 67456
        325: data_ff <= 24'hFF53D9; // -44071
        326: data_ff <= 24'h006D9B; // 28059
        327: data_ff <= 24'hFFBCDE; // -17186
        328: data_ff <= 24'h002718; // 10008
        329: data_ff <= 24'hFFEAA2; // -5470
        330: data_ff <= 24'h000ACB; // 2763
        331: data_ff <= 24'hFFFB12; // -1262
        332: data_ff <= 24'h0001F8; // 504
        333: data_ff <= 24'hFFFF5C; // -164
        334: data_ff <= 24'h000024; // 36
        335: data_ff <= 24'hFFFFFE; // -2
        336: data_ff <= 24'h099CC3; // 629955
        337: data_ff <= 24'hFBBD5B; // -279205
        338: data_ff <= 24'h0287D7; // 165847
        339: data_ff <= 24'hFE5DFE; // -107010
        340: data_ff <= 24'h01133D; // 70461
        341: data_ff <= 24'hFF4C4B; // -46005
        342: data_ff <= 24'h00725C; // 29276
        343: data_ff <= 24'hFFB9FC; // -17924
        344: data_ff <= 24'h0028C2; // 10434
        345: data_ff <= 24'hFFE9BA; // -5702
        346: data_ff <= 24'h000B40; // 2880
        347: data_ff <= 24'hFFFADD; // -1315
        348: data_ff <= 24'h00020D; // 525
        349: data_ff <= 24'hFFFF54; // -172
        350: data_ff <= 24'h000026; // 38
        351: data_ff <= 24'hFFFFFE; // -2
        352: data_ff <= 24'h0A1926; // 661798
        353: data_ff <= 24'hFB8B3A; // -292038
        354: data_ff <= 24'h02A484; // 173188
        355: data_ff <= 24'hFE4BEC; // -111636
        356: data_ff <= 24'h011EEE; // 73454
        357: data_ff <= 24'hFF44C4; // -47932
        358: data_ff <= 24'h007718; // 30488
        359: data_ff <= 24'hFFB71D; // -18659
        360: data_ff <= 24'h002A6B; // 10859
        361: data_ff <= 24'hFFE8D2; // -5934
        362: data_ff <= 24'h000BB4; // 2996
        363: data_ff <= 24'hFFFAA7; // -1369
        364: data_ff <= 24'h000223; // 547
        365: data_ff <= 24'hFFFF4D; // -179
        366: data_ff <= 24'h000027; // 39
        367: data_ff <= 24'hFFFFFD; // -3
        368: data_ff <= 24'h0A9668; // 693864
        369: data_ff <= 24'hFB5926; // -304858
        370: data_ff <= 24'h02C11A; // 180506
        371: data_ff <= 24'hFE39EB; // -116245
        372: data_ff <= 24'h012A93; // 76435
        373: data_ff <= 24'hFF3D44; // -49852
        374: data_ff <= 24'h007BD0; // 31696
        375: data_ff <= 24'hFFB440; // -19392
        376: data_ff <= 24'h002C13; // 11283
        377: data_ff <= 24'hFFE7EC; // -6164
        378: data_ff <= 24'h000C29; // 3113
        379: data_ff <= 24'hFFFA72; // -1422
        380: data_ff <= 24'h000239; // 569
        381: data_ff <= 24'hFFFF46; // -186
        382: data_ff <= 24'h000029; // 41
        383: data_ff <= 24'hFFFFFD; // -3
        384: data_ff <= 24'h0B1483; // 726147
        385: data_ff <= 24'hFB2725; // -317659
        386: data_ff <= 24'h02DD95; // 187797
        387: data_ff <= 24'hFE2800; // -120832
        388: data_ff <= 24'h01362A; // 79402
        389: data_ff <= 24'hFF35CE; // -51762
        390: data_ff <= 24'h008082; // 32898
        391: data_ff <= 24'hFFB166; // -20122
        392: data_ff <= 24'h002DBA; // 11706
        393: data_ff <= 24'hFFE705; // -6395
        394: data_ff <= 24'h000C9D; // 3229
        395: data_ff <= 24'hFFFA3C; // -1476
        396: data_ff <= 24'h00024E; // 590
        397: data_ff <= 24'hFFFF3E; // -194
        398: data_ff <= 24'h00002B; // 43
        399: data_ff <= 24'hFFFFFD; // -3
        400: data_ff <= 24'h0B9370; // 758640
        401: data_ff <= 24'hFAF53D; // -330435
        402: data_ff <= 24'h02F9F3; // 195059
        403: data_ff <= 24'hFE162A; // -125398
        404: data_ff <= 24'h0141B2; // 82354
        405: data_ff <= 24'hFF2E61; // -53663
        406: data_ff <= 24'h00852F; // 34095
        407: data_ff <= 24'hFFAE8F; // -20849
        408: data_ff <= 24'h002F5F; // 12127
        409: data_ff <= 24'hFFE620; // -6624
        410: data_ff <= 24'h000D11; // 3345
        411: data_ff <= 24'hFFFA07; // -1529
        412: data_ff <= 24'h000264; // 612
        413: data_ff <= 24'hFFFF37; // -201
        414: data_ff <= 24'h00002D; // 45
        415: data_ff <= 24'hFFFFFD; // -3
        416: data_ff <= 24'h0C132B; // 791339
        417: data_ff <= 24'hFAC371; // -343183
        418: data_ff <= 24'h031630; // 202288
        419: data_ff <= 24'hFE046C; // -129940
        420: data_ff <= 24'h014D2A; // 85290
        421: data_ff <= 24'hFF26FF; // -55553
        422: data_ff <= 24'h0089D5; // 35285
        423: data_ff <= 24'hFFABBC; // -21572
        424: data_ff <= 24'h003102; // 12546
        425: data_ff <= 24'hFFE53B; // -6853
        426: data_ff <= 24'h000D85; // 3461
        427: data_ff <= 24'hFFF9D2; // -1582
        428: data_ff <= 24'h00027A; // 634
        429: data_ff <= 24'hFFFF30; // -208
        430: data_ff <= 24'h00002E; // 46
        431: data_ff <= 24'hFFFFFD; // -3
        432: data_ff <= 24'h0C93AC; // 824236
        433: data_ff <= 24'hFA91C6; // -355898
        434: data_ff <= 24'h03324A; // 209482
        435: data_ff <= 24'hFDF2C9; // -134455
        436: data_ff <= 24'h015890; // 88208
        437: data_ff <= 24'hFF1FA8; // -57432
        438: data_ff <= 24'h008E75; // 36469
        439: data_ff <= 24'hFFA8EC; // -22292
        440: data_ff <= 24'h0032A3; // 12963
        441: data_ff <= 24'hFFE457; // -7081
        442: data_ff <= 24'h000DF9; // 3577
        443: data_ff <= 24'hFFF99C; // -1636
        444: data_ff <= 24'h00028F; // 655
        445: data_ff <= 24'hFFFF28; // -216
        446: data_ff <= 24'h000030; // 48
        447: data_ff <= 24'hFFFFFD; // -3
        448: data_ff <= 24'h0D14ED; // 857325
        449: data_ff <= 24'hFA6043; // -368573
        450: data_ff <= 24'h034E3E; // 216638
        451: data_ff <= 24'hFDE141; // -138943
        452: data_ff <= 24'h0163E3; // 91107
        453: data_ff <= 24'hFF185C; // -59300
        454: data_ff <= 24'h00930D; // 37645
        455: data_ff <= 24'hFFA621; // -23007
        456: data_ff <= 24'h003442; // 13378
        457: data_ff <= 24'hFFE375; // -7307
        458: data_ff <= 24'h000E6C; // 3692
        459: data_ff <= 24'hFFF967; // -1689
        460: data_ff <= 24'h0002A5; // 677
        461: data_ff <= 24'hFFFF21; // -223
        462: data_ff <= 24'h000032; // 50
        463: data_ff <= 24'hFFFFFC; // -4
        464: data_ff <= 24'h0D96EA; // 890602
        465: data_ff <= 24'hFA2EEB; // -381205
        466: data_ff <= 24'h036A07; // 223751
        467: data_ff <= 24'hFDCFD7; // -143401
        468: data_ff <= 24'h016F22; // 93986
        469: data_ff <= 24'hFF111E; // -61154
        470: data_ff <= 24'h00979E; // 38814
        471: data_ff <= 24'hFFA35A; // -23718
        472: data_ff <= 24'h0035DE; // 13790
        473: data_ff <= 24'hFFE293; // -7533
        474: data_ff <= 24'h000EDE; // 3806
        475: data_ff <= 24'hFFF932; // -1742
        476: data_ff <= 24'h0002BB; // 699
        477: data_ff <= 24'hFFFF19; // -231
        478: data_ff <= 24'h000034; // 52
        479: data_ff <= 24'hFFFFFC; // -4
        480: data_ff <= 24'h0E199A; // 924058
        481: data_ff <= 24'hF9FDC4; // -393788
        482: data_ff <= 24'h0385A5; // 230821
        483: data_ff <= 24'hFDBE8D; // -147827
        484: data_ff <= 24'h017A4C; // 96844
        485: data_ff <= 24'hFF09ED; // -62995
        486: data_ff <= 24'h009C26; // 39974
        487: data_ff <= 24'hFFA098; // -24424
        488: data_ff <= 24'h003778; // 14200
        489: data_ff <= 24'hFFE1B3; // -7757
        490: data_ff <= 24'h000F51; // 3921
        491: data_ff <= 24'hFFF8FD; // -1795
        492: data_ff <= 24'h0002D0; // 720
        493: data_ff <= 24'hFFFF12; // -238
        494: data_ff <= 24'h000036; // 54
        495: data_ff <= 24'hFFFFFC; // -4
        496: data_ff <= 24'h0E9CF8; // 957688
        497: data_ff <= 24'hF9CCD3; // -406317
        498: data_ff <= 24'h03A113; // 237843
        499: data_ff <= 24'hFDAD65; // -152219
        500: data_ff <= 24'h018560; // 99680
        501: data_ff <= 24'hFF02CB; // -64821
        502: data_ff <= 24'h00A0A6; // 41126
        503: data_ff <= 24'hFF9DDB; // -25125
        504: data_ff <= 24'h003910; // 14608
        505: data_ff <= 24'hFFE0D3; // -7981
        506: data_ff <= 24'h000FC2; // 4034
        507: data_ff <= 24'hFFF8C9; // -1847
        508: data_ff <= 24'h0002E6; // 742
        509: data_ff <= 24'hFFFF0B; // -245
        510: data_ff <= 24'h000038; // 56
        511: data_ff <= 24'hFFFFFC; // -4
        512: data_ff <= 24'h0F20FD; // 991485
        513: data_ff <= 24'hF99C1C; // -418788
        514: data_ff <= 24'h03BC4F; // 244815
        515: data_ff <= 24'hFD9C60; // -156576
        516: data_ff <= 24'h01905C; // 102492
        517: data_ff <= 24'hFEFBB8; // -66632
        518: data_ff <= 24'h00A51C; // 42268
        519: data_ff <= 24'hFF9B23; // -25821
        520: data_ff <= 24'h003AA4; // 15012
        521: data_ff <= 24'hFFDFF6; // -8202
        522: data_ff <= 24'h001033; // 4147
        523: data_ff <= 24'hFFF894; // -1900
        524: data_ff <= 24'h0002FB; // 763
        525: data_ff <= 24'hFFFF03; // -253
        526: data_ff <= 24'h00003A; // 58
        527: data_ff <= 24'hFFFFFC; // -4
        528: data_ff <= 24'h0FA5A3; // 1025443
        529: data_ff <= 24'hF96BA6; // -431194
        530: data_ff <= 24'h03D755; // 251733
        531: data_ff <= 24'hFD8B80; // -160896
        532: data_ff <= 24'h019B3E; // 105278
        533: data_ff <= 24'hFEF4B5; // -68427
        534: data_ff <= 24'h00A988; // 43400
        535: data_ff <= 24'hFF9871; // -26511
        536: data_ff <= 24'h003C36; // 15414
        537: data_ff <= 24'hFFDF19; // -8423
        538: data_ff <= 24'h0010A3; // 4259
        539: data_ff <= 24'hFFF860; // -1952
        540: data_ff <= 24'h000311; // 785
        541: data_ff <= 24'hFFFEFC; // -260
        542: data_ff <= 24'h00003C; // 60
        543: data_ff <= 24'hFFFFFC; // -4
        544: data_ff <= 24'h102AE3; // 1059555
        545: data_ff <= 24'hF93B75; // -443531
        546: data_ff <= 24'h03F223; // 258595
        547: data_ff <= 24'hFD7AC8; // -165176
        548: data_ff <= 24'h01A607; // 108039
        549: data_ff <= 24'hFEEDC3; // -70205
        550: data_ff <= 24'h00ADEA; // 44522
        551: data_ff <= 24'hFF95C5; // -27195
        552: data_ff <= 24'h003DC4; // 15812
        553: data_ff <= 24'hFFDE3F; // -8641
        554: data_ff <= 24'h001113; // 4371
        555: data_ff <= 24'hFFF82C; // -2004
        556: data_ff <= 24'h000326; // 806
        557: data_ff <= 24'hFFFEF4; // -268
        558: data_ff <= 24'h00003D; // 61
        559: data_ff <= 24'hFFFFFB; // -5
        560: data_ff <= 24'h10B0B6; // 1093814
        561: data_ff <= 24'hF90B8D; // -455795
        562: data_ff <= 24'h040CB6; // 265398
        563: data_ff <= 24'hFD6A38; // -169416
        564: data_ff <= 24'h01B0B4; // 110772
        565: data_ff <= 24'hFEE6E2; // -71966
        566: data_ff <= 24'h00B241; // 45633
        567: data_ff <= 24'hFF931F; // -27873
        568: data_ff <= 24'h003F4F; // 16207
        569: data_ff <= 24'hFFDD66; // -8858
        570: data_ff <= 24'h001182; // 4482
        571: data_ff <= 24'hFFF7F8; // -2056
        572: data_ff <= 24'h00033C; // 828
        573: data_ff <= 24'hFFFEED; // -275
        574: data_ff <= 24'h00003F; // 63
        575: data_ff <= 24'hFFFFFB; // -5
        576: data_ff <= 24'h113717; // 1128215
        577: data_ff <= 24'hF8DBF6; // -467978
        578: data_ff <= 24'h04270A; // 272138
        579: data_ff <= 24'hFD59D4; // -173612
        580: data_ff <= 24'h01BB45; // 113477
        581: data_ff <= 24'hFEE014; // -73708
        582: data_ff <= 24'h00B68D; // 46733
        583: data_ff <= 24'hFF9080; // -28544
        584: data_ff <= 24'h0040D6; // 16598
        585: data_ff <= 24'hFFDC8F; // -9073
        586: data_ff <= 24'h0011F0; // 4592
        587: data_ff <= 24'hFFF7C5; // -2107
        588: data_ff <= 24'h000351; // 849
        589: data_ff <= 24'hFFFEE5; // -283
        590: data_ff <= 24'h000041; // 65
        591: data_ff <= 24'hFFFFFB; // -5
        592: data_ff <= 24'h11BDFE; // 1162750
        593: data_ff <= 24'hF8ACB2; // -480078
        594: data_ff <= 24'h04411D; // 278813
        595: data_ff <= 24'hFD499D; // -177763
        596: data_ff <= 24'h01C5B7; // 116151
        597: data_ff <= 24'hFED959; // -75431
        598: data_ff <= 24'h00BACD; // 47821
        599: data_ff <= 24'hFF8DE8; // -29208
        600: data_ff <= 24'h004259; // 16985
        601: data_ff <= 24'hFFDBBA; // -9286
        602: data_ff <= 24'h00125D; // 4701
        603: data_ff <= 24'hFFF792; // -2158
        604: data_ff <= 24'h000366; // 870
        605: data_ff <= 24'hFFFEDE; // -290
        606: data_ff <= 24'h000043; // 67
        607: data_ff <= 24'hFFFFFB; // -5
        608: data_ff <= 24'h124563; // 1197411
        609: data_ff <= 24'hF87DC8; // -492088
        610: data_ff <= 24'h045AEC; // 285420
        611: data_ff <= 24'hFD3995; // -181867
        612: data_ff <= 24'h01D00B; // 118795
        613: data_ff <= 24'hFED2B2; // -77134
        614: data_ff <= 24'h00BF01; // 48897
        615: data_ff <= 24'hFF8B57; // -29865
        616: data_ff <= 24'h0043D8; // 17368
        617: data_ff <= 24'hFFDAE7; // -9497
        618: data_ff <= 24'h0012C9; // 4809
        619: data_ff <= 24'hFFF75F; // -2209
        620: data_ff <= 24'h00037B; // 891
        621: data_ff <= 24'hFFFED7; // -297
        622: data_ff <= 24'h000045; // 69
        623: data_ff <= 24'hFFFFFB; // -5
        624: data_ff <= 24'h12CD42; // 1232194
        625: data_ff <= 24'hF84F3D; // -504003
        626: data_ff <= 24'h047474; // 291956
        627: data_ff <= 24'hFD29BD; // -185923
        628: data_ff <= 24'h01DA3E; // 121406
        629: data_ff <= 24'hFECC20; // -78816
        630: data_ff <= 24'h00C327; // 49959
        631: data_ff <= 24'hFF88CE; // -30514
        632: data_ff <= 24'h004553; // 17747
        633: data_ff <= 24'hFFDA16; // -9706
        634: data_ff <= 24'h001334; // 4916
        635: data_ff <= 24'hFFF72D; // -2259
        636: data_ff <= 24'h000390; // 912
        637: data_ff <= 24'hFFFECF; // -305
        638: data_ff <= 24'h000047; // 71
        639: data_ff <= 24'hFFFFFA; // -6
        640: data_ff <= 24'h135592; // 1267090
        641: data_ff <= 24'hF82116; // -515818
        642: data_ff <= 24'h048DB1; // 298417
        643: data_ff <= 24'hFD1A17; // -189929
        644: data_ff <= 24'h01E450; // 123984
        645: data_ff <= 24'hFEC5A3; // -80477
        646: data_ff <= 24'h00C741; // 51009
        647: data_ff <= 24'hFF864D; // -31155
        648: data_ff <= 24'h0046CA; // 18122
        649: data_ff <= 24'hFFD947; // -9913
        650: data_ff <= 24'h00139E; // 5022
        651: data_ff <= 24'hFFF6FB; // -2309
        652: data_ff <= 24'h0003A5; // 933
        653: data_ff <= 24'hFFFEC8; // -312
        654: data_ff <= 24'h000049; // 73
        655: data_ff <= 24'hFFFFFA; // -6
        656: data_ff <= 24'h13DE4C; // 1302092
        657: data_ff <= 24'hF7F358; // -527528
        658: data_ff <= 24'h04A6A2; // 304802
        659: data_ff <= 24'hFD0AA6; // -193882
        660: data_ff <= 24'h01EE3F; // 126527
        661: data_ff <= 24'hFEBF3D; // -82115
        662: data_ff <= 24'h00CB4C; // 52044
        663: data_ff <= 24'hFF83D3; // -31789
        664: data_ff <= 24'h00483C; // 18492
        665: data_ff <= 24'hFFD87B; // -10117
        666: data_ff <= 24'h001408; // 5128
        667: data_ff <= 24'hFFF6CA; // -2358
        668: data_ff <= 24'h0003B9; // 953
        669: data_ff <= 24'hFFFEC1; // -319
        670: data_ff <= 24'h00004B; // 75
        671: data_ff <= 24'hFFFFFA; // -6
        672: data_ff <= 24'h14676A; // 1337194
        673: data_ff <= 24'hF7C608; // -539128
        674: data_ff <= 24'h04BF42; // 311106
        675: data_ff <= 24'hFCFB6C; // -197780
        676: data_ff <= 24'h01F80A; // 129034
        677: data_ff <= 24'hFEB8EE; // -83730
        678: data_ff <= 24'h00CF49; // 53065
        679: data_ff <= 24'hFF8163; // -32413
        680: data_ff <= 24'h0049AA; // 18858
        681: data_ff <= 24'hFFD7B1; // -10319
        682: data_ff <= 24'h00146F; // 5231
        683: data_ff <= 24'hFFF699; // -2407
        684: data_ff <= 24'h0003CE; // 974
        685: data_ff <= 24'hFFFEB9; // -327
        686: data_ff <= 24'h00004D; // 77
        687: data_ff <= 24'hFFFFFA; // -6
        688: data_ff <= 24'h14F0E4; // 1372388
        689: data_ff <= 24'hF7992C; // -550612
        690: data_ff <= 24'h04D78F; // 317327
        691: data_ff <= 24'hFCEC69; // -201623
        692: data_ff <= 24'h0201B0; // 131504
        693: data_ff <= 24'hFEB2B7; // -85321
        694: data_ff <= 24'h00D337; // 54071
        695: data_ff <= 24'hFF7EFB; // -33029
        696: data_ff <= 24'h004B12; // 19218
        697: data_ff <= 24'hFFD6E9; // -10519
        698: data_ff <= 24'h0014D6; // 5334
        699: data_ff <= 24'hFFF669; // -2455
        700: data_ff <= 24'h0003E2; // 994
        701: data_ff <= 24'hFFFEB2; // -334
        702: data_ff <= 24'h00004F; // 79
        703: data_ff <= 24'hFFFFFA; // -6
        704: data_ff <= 24'h157AB4; // 1407668
        705: data_ff <= 24'hF76CC8; // -561976
        706: data_ff <= 24'h04EF87; // 323463
        707: data_ff <= 24'hFCDDA0; // -205408
        708: data_ff <= 24'h020B30; // 133936
        709: data_ff <= 24'hFEAC98; // -86888
        710: data_ff <= 24'h00D716; // 55062
        711: data_ff <= 24'hFF7C9C; // -33636
        712: data_ff <= 24'h004C75; // 19573
        713: data_ff <= 24'hFFD624; // -10716
        714: data_ff <= 24'h00153C; // 5436
        715: data_ff <= 24'hFFF639; // -2503
        716: data_ff <= 24'h0003F6; // 1014
        717: data_ff <= 24'hFFFEAB; // -341
        718: data_ff <= 24'h000051; // 81
        719: data_ff <= 24'hFFFFF9; // -7
        720: data_ff <= 24'h1604D2; // 1443026
        721: data_ff <= 24'hF740E2; // -573214
        722: data_ff <= 24'h050726; // 329510
        723: data_ff <= 24'hFCCF12; // -209134
        724: data_ff <= 24'h021488; // 136328
        725: data_ff <= 24'hFEA693; // -88429
        726: data_ff <= 24'h00DAE5; // 56037
        727: data_ff <= 24'hFF7A47; // -34233
        728: data_ff <= 24'h004DD4; // 19924
        729: data_ff <= 24'hFFD562; // -10910
        730: data_ff <= 24'h0015A0; // 5536
        731: data_ff <= 24'hFFF609; // -2551
        732: data_ff <= 24'h00040A; // 1034
        733: data_ff <= 24'hFFFEA4; // -348
        734: data_ff <= 24'h000053; // 83
        735: data_ff <= 24'hFFFFF9; // -7
        736: data_ff <= 24'h168F37; // 1478455
        737: data_ff <= 24'hF7157F; // -584321
        738: data_ff <= 24'h051E69; // 335465
        739: data_ff <= 24'hFCC0C2; // -212798
        740: data_ff <= 24'h021DB8; // 138680
        741: data_ff <= 24'hFEA0A8; // -89944
        742: data_ff <= 24'h00DEA4; // 56996
        743: data_ff <= 24'hFF77FB; // -34821
        744: data_ff <= 24'h004F2C; // 20268
        745: data_ff <= 24'hFFD4A3; // -11101
        746: data_ff <= 24'h001603; // 5635
        747: data_ff <= 24'hFFF5DB; // -2597
        748: data_ff <= 24'h00041E; // 1054
        749: data_ff <= 24'hFFFE9D; // -355
        750: data_ff <= 24'h000055; // 85
        751: data_ff <= 24'hFFFFF9; // -7
        752: data_ff <= 24'h1719DB; // 1513947
        753: data_ff <= 24'hF6EAA4; // -595292
        754: data_ff <= 24'h05354E; // 341326
        755: data_ff <= 24'hFCB2B1; // -216399
        756: data_ff <= 24'h0226BF; // 140991
        757: data_ff <= 24'hFE9AD8; // -91432
        758: data_ff <= 24'h00E252; // 57938
        759: data_ff <= 24'hFF75B9; // -35399
        760: data_ff <= 24'h00507F; // 20607
        761: data_ff <= 24'hFFD3E7; // -11289
        762: data_ff <= 24'h001664; // 5732
        763: data_ff <= 24'hFFF5AC; // -2644
        764: data_ff <= 24'h000432; // 1074
        765: data_ff <= 24'hFFFE95; // -363
        766: data_ff <= 24'h000057; // 87
        767: data_ff <= 24'hFFFFF9; // -7
        768: data_ff <= 24'h17A4B8; // 1549496
        769: data_ff <= 24'hF6C057; // -606121
        770: data_ff <= 24'h054BD2; // 347090
        771: data_ff <= 24'hFCA4E1; // -219935
        772: data_ff <= 24'h022F9A; // 143258
        773: data_ff <= 24'hFE9524; // -92892
        774: data_ff <= 24'h00E5EF; // 58863
        775: data_ff <= 24'hFF7382; // -35966
        776: data_ff <= 24'h0051CD; // 20941
        777: data_ff <= 24'hFFD32E; // -11474
        778: data_ff <= 24'h0016C4; // 5828
        779: data_ff <= 24'hFFF57F; // -2689
        780: data_ff <= 24'h000445; // 1093
        781: data_ff <= 24'hFFFE8E; // -370
        782: data_ff <= 24'h000059; // 89
        783: data_ff <= 24'hFFFFF8; // -8
        784: data_ff <= 24'h182FC6; // 1585094
        785: data_ff <= 24'hF6969C; // -616804
        786: data_ff <= 24'h0561F2; // 352754
        787: data_ff <= 24'hFC9753; // -223405
        788: data_ff <= 24'h02384A; // 145482
        789: data_ff <= 24'hFE8F8C; // -94324
        790: data_ff <= 24'h00E97A; // 59770
        791: data_ff <= 24'hFF7155; // -36523
        792: data_ff <= 24'h005314; // 21268
        793: data_ff <= 24'hFFD278; // -11656
        794: data_ff <= 24'h001723; // 5923
        795: data_ff <= 24'hFFF552; // -2734
        796: data_ff <= 24'h000458; // 1112
        797: data_ff <= 24'hFFFE88; // -376
        798: data_ff <= 24'h00005B; // 91
        799: data_ff <= 24'hFFFFF8; // -8
        800: data_ff <= 24'h18BAFE; // 1620734
        801: data_ff <= 24'hF66D78; // -627336
        802: data_ff <= 24'h0577AB; // 358315
        803: data_ff <= 24'hFC8A09; // -226807
        804: data_ff <= 24'h0240CC; // 147660
        805: data_ff <= 24'hFE8A11; // -95727
        806: data_ff <= 24'h00ECF2; // 60658
        807: data_ff <= 24'hFF6F33; // -37069
        808: data_ff <= 24'h005455; // 21589
        809: data_ff <= 24'hFFD1C5; // -11835
        810: data_ff <= 24'h001780; // 6016
        811: data_ff <= 24'hFFF526; // -2778
        812: data_ff <= 24'h00046B; // 1131
        813: data_ff <= 24'hFFFE81; // -383
        814: data_ff <= 24'h00005D; // 93
        815: data_ff <= 24'hFFFFF8; // -8
        816: data_ff <= 24'h194658; // 1656408
        817: data_ff <= 24'hF644F2; // -637710
        818: data_ff <= 24'h058CFA; // 363770
        819: data_ff <= 24'hFC7D06; // -230138
        820: data_ff <= 24'h024920; // 149792
        821: data_ff <= 24'hFE84B4; // -97100
        822: data_ff <= 24'h00F059; // 61529
        823: data_ff <= 24'hFF6D1D; // -37603
        824: data_ff <= 24'h005590; // 21904
        825: data_ff <= 24'hFFD116; // -12010
        826: data_ff <= 24'h0017DB; // 6107
        827: data_ff <= 24'hFFF4FA; // -2822
        828: data_ff <= 24'h00047E; // 1150
        829: data_ff <= 24'hFFFE7A; // -390
        830: data_ff <= 24'h00005F; // 95
        831: data_ff <= 24'hFFFFF8; // -8
        832: data_ff <= 24'h19D1CD; // 1692109
        833: data_ff <= 24'hF61D0D; // -647923
        834: data_ff <= 24'h05A1DD; // 369117
        835: data_ff <= 24'hFC704A; // -233398
        836: data_ff <= 24'h025146; // 151878
        837: data_ff <= 24'hFE7F75; // -98443
        838: data_ff <= 24'h00F3AB; // 62379
        839: data_ff <= 24'hFF6B12; // -38126
        840: data_ff <= 24'h0056C4; // 22212
        841: data_ff <= 24'hFFD06A; // -12182
        842: data_ff <= 24'h001835; // 6197
        843: data_ff <= 24'hFFF4CF; // -2865
        844: data_ff <= 24'h000490; // 1168
        845: data_ff <= 24'hFFFE73; // -397
        846: data_ff <= 24'h000060; // 96
        847: data_ff <= 24'hFFFFF7; // -9
        848: data_ff <= 24'h1A5D56; // 1727830
        849: data_ff <= 24'hF5F5CF; // -657969
        850: data_ff <= 24'h05B650; // 374352
        851: data_ff <= 24'hFC63D8; // -236584
        852: data_ff <= 24'h02593A; // 153914
        853: data_ff <= 24'hFE7A56; // -99754
        854: data_ff <= 24'h00F6EB; // 63211
        855: data_ff <= 24'hFF6912; // -38638
        856: data_ff <= 24'h0057F2; // 22514
        857: data_ff <= 24'hFFCFC1; // -12351
        858: data_ff <= 24'h00188C; // 6284
        859: data_ff <= 24'hFFF4A5; // -2907
        860: data_ff <= 24'h0004A2; // 1186
        861: data_ff <= 24'hFFFE6D; // -403
        862: data_ff <= 24'h000062; // 98
        863: data_ff <= 24'hFFFFF7; // -9
        864: data_ff <= 24'h1AE8EA; // 1763562
        865: data_ff <= 24'hF5CF3D; // -667843
        866: data_ff <= 24'h05CA52; // 379474
        867: data_ff <= 24'hFC57B1; // -239695
        868: data_ff <= 24'h0260FE; // 155902
        869: data_ff <= 24'hFE7557; // -101033
        870: data_ff <= 24'h00FA16; // 64022
        871: data_ff <= 24'hFF671F; // -39137
        872: data_ff <= 24'h005918; // 22808
        873: data_ff <= 24'hFFCF1C; // -12516
        874: data_ff <= 24'h0018E3; // 6371
        875: data_ff <= 24'hFFF47C; // -2948
        876: data_ff <= 24'h0004B4; // 1204
        877: data_ff <= 24'hFFFE66; // -410
        878: data_ff <= 24'h000064; // 100
        879: data_ff <= 24'hFFFFF7; // -9
        880: data_ff <= 24'h1B7484; // 1799300
        881: data_ff <= 24'hF5A95D; // -677539
        882: data_ff <= 24'h05DDE0; // 384480
        883: data_ff <= 24'hFC4BD6; // -242730
        884: data_ff <= 24'h02688F; // 157839
        885: data_ff <= 24'hFE7078; // -102280
        886: data_ff <= 24'h00FD2D; // 64813
        887: data_ff <= 24'hFF6538; // -39624
        888: data_ff <= 24'h005A38; // 23096
        889: data_ff <= 24'hFFCE7B; // -12677
        890: data_ff <= 24'h001937; // 6455
        891: data_ff <= 24'hFFF453; // -2989
        892: data_ff <= 24'h0004C5; // 1221
        893: data_ff <= 24'hFFFE5F; // -417
        894: data_ff <= 24'h000066; // 102
        895: data_ff <= 24'hFFFFF7; // -9
        896: data_ff <= 24'h1C001A; // 1835034
        897: data_ff <= 24'hF58433; // -687053
        898: data_ff <= 24'h05F0F6; // 389366
        899: data_ff <= 24'hFC404A; // -245686
        900: data_ff <= 24'h026FED; // 159725
        901: data_ff <= 24'hFE6BBA; // -103494
        902: data_ff <= 24'h01002F; // 65583
        903: data_ff <= 24'hFF635D; // -40099
        904: data_ff <= 24'h005B51; // 23377
        905: data_ff <= 24'hFFCDDE; // -12834
        906: data_ff <= 24'h001989; // 6537
        907: data_ff <= 24'hFFF42B; // -3029
        908: data_ff <= 24'h0004D6; // 1238
        909: data_ff <= 24'hFFFE59; // -423
        910: data_ff <= 24'h000068; // 104
        911: data_ff <= 24'hFFFFF6; // -10
        912: data_ff <= 24'h1C8BA5; // 1870757
        913: data_ff <= 24'hF55FC3; // -696381
        914: data_ff <= 24'h060393; // 394131
        915: data_ff <= 24'hFC350D; // -248563
        916: data_ff <= 24'h027716; // 161558
        917: data_ff <= 24'hFE671F; // -104673
        918: data_ff <= 24'h01031C; // 66332
        919: data_ff <= 24'hFF618F; // -40561
        920: data_ff <= 24'h005C62; // 23650
        921: data_ff <= 24'hFFCD45; // -12987
        922: data_ff <= 24'h0019DA; // 6618
        923: data_ff <= 24'hFFF405; // -3067
        924: data_ff <= 24'h0004E7; // 1255
        925: data_ff <= 24'hFFFE53; // -429
        926: data_ff <= 24'h00006A; // 106
        927: data_ff <= 24'hFFFFF6; // -10
        928: data_ff <= 24'h1D171E; // 1906462
        929: data_ff <= 24'hF53C14; // -705516
        930: data_ff <= 24'h0615B3; // 398771
        931: data_ff <= 24'hFC2A22; // -251358
        932: data_ff <= 24'h027E0A; // 163338
        933: data_ff <= 24'hFE62A6; // -105818
        934: data_ff <= 24'h0105F3; // 67059
        935: data_ff <= 24'hFF5FCF; // -41009
        936: data_ff <= 24'h005D6B; // 23915
        937: data_ff <= 24'hFFCCB0; // -13136
        938: data_ff <= 24'h001A28; // 6696
        939: data_ff <= 24'hFFF3DF; // -3105
        940: data_ff <= 24'h0004F8; // 1272
        941: data_ff <= 24'hFFFE4D; // -435
        942: data_ff <= 24'h00006C; // 108
        943: data_ff <= 24'hFFFFF6; // -10
        944: data_ff <= 24'h1DA27E; // 1942142
        945: data_ff <= 24'hF5192B; // -714453
        946: data_ff <= 24'h062755; // 403285
        947: data_ff <= 24'hFC1F89; // -254071
        948: data_ff <= 24'h0284C7; // 165063
        949: data_ff <= 24'hFE5E50; // -106928
        950: data_ff <= 24'h0108B4; // 67764
        951: data_ff <= 24'hFF5E1C; // -41444
        952: data_ff <= 24'h005E6D; // 24173
        953: data_ff <= 24'hFFCC1F; // -13281
        954: data_ff <= 24'h001A75; // 6773
        955: data_ff <= 24'hFFF3BA; // -3142
        956: data_ff <= 24'h000508; // 1288
        957: data_ff <= 24'hFFFE47; // -441
        958: data_ff <= 24'h00006E; // 110
        959: data_ff <= 24'hFFFFF5; // -11
        960: data_ff <= 24'h1E2DBC; // 1977788
        961: data_ff <= 24'hF4F70B; // -723189
        962: data_ff <= 24'h063875; // 407669
        963: data_ff <= 24'hFC1545; // -256699
        964: data_ff <= 24'h028B4D; // 166733
        965: data_ff <= 24'hFE5A1E; // -108002
        966: data_ff <= 24'h010B5E; // 68446
        967: data_ff <= 24'hFF5C76; // -41866
        968: data_ff <= 24'h005F68; // 24424
        969: data_ff <= 24'hFFCB92; // -13422
        970: data_ff <= 24'h001ABF; // 6847
        971: data_ff <= 24'hFFF395; // -3179
        972: data_ff <= 24'h000518; // 1304
        973: data_ff <= 24'hFFFE41; // -447
        974: data_ff <= 24'h00006F; // 111
        975: data_ff <= 24'hFFFFF5; // -11
        976: data_ff <= 24'h1EB8D2; // 2013394
        977: data_ff <= 24'hF4D5BB; // -731717
        978: data_ff <= 24'h064911; // 411921
        979: data_ff <= 24'hFC0B57; // -259241
        980: data_ff <= 24'h02919A; // 168346
        981: data_ff <= 24'hFE5611; // -109039
        982: data_ff <= 24'h010DF1; // 69105
        983: data_ff <= 24'hFF5ADF; // -42273
        984: data_ff <= 24'h00605A; // 24666
        985: data_ff <= 24'hFFCB09; // -13559
        986: data_ff <= 24'h001B07; // 6919
        987: data_ff <= 24'hFFF372; // -3214
        988: data_ff <= 24'h000527; // 1319
        989: data_ff <= 24'hFFFE3B; // -453
        990: data_ff <= 24'h000071; // 113
        991: data_ff <= 24'hFFFFF5; // -11
        992: data_ff <= 24'h1F43B6; // 2048950
        993: data_ff <= 24'hF4B53F; // -740033
        994: data_ff <= 24'h065927; // 416039
        995: data_ff <= 24'hFC01C1; // -261695
        996: data_ff <= 24'h0297AE; // 169902
        997: data_ff <= 24'hFE5229; // -110039
        998: data_ff <= 24'h01106D; // 69741
        999: data_ff <= 24'hFF5955; // -42667
        1000: data_ff <= 24'h006144; // 24900
        1001: data_ff <= 24'hFFCA85; // -13691
        1002: data_ff <= 24'h001B4D; // 6989
        1003: data_ff <= 24'hFFF350; // -3248
        1004: data_ff <= 24'h000536; // 1334
        1005: data_ff <= 24'hFFFE35; // -459
        1006: data_ff <= 24'h000073; // 115
        1007: data_ff <= 24'hFFFFF5; // -11
        1008: data_ff <= 24'h1FCE63; // 2084451
        1009: data_ff <= 24'hF4959B; // -748133
        1010: data_ff <= 24'h0668B5; // 420021
        1011: data_ff <= 24'hFBF883; // -264061
        1012: data_ff <= 24'h029D88; // 171400
        1013: data_ff <= 24'hFE4E66; // -111002
        1014: data_ff <= 24'h0112D1; // 70353
        1015: data_ff <= 24'hFF57DA; // -43046
        1016: data_ff <= 24'h006225; // 25125
        1017: data_ff <= 24'hFFCA05; // -13819
        1018: data_ff <= 24'h001B91; // 7057
        1019: data_ff <= 24'hFFF32F; // -3281
        1020: data_ff <= 24'h000545; // 1349
        1021: data_ff <= 24'hFFFE2F; // -465
        1022: data_ff <= 24'h000075; // 117
        1023: data_ff <= 24'hFFFFF4; // -12
        1024: data_ff <= 24'h2058CF; // 2119887
        1025: data_ff <= 24'hF476D5; // -756011
        1026: data_ff <= 24'h0677B7; // 423863
        1027: data_ff <= 24'hFBEF9F; // -266337
        1028: data_ff <= 24'h02A327; // 172839
        1029: data_ff <= 24'hFE4ACA; // -111926
        1030: data_ff <= 24'h01151D; // 70941
        1031: data_ff <= 24'hFF566E; // -43410
        1032: data_ff <= 24'h0062FF; // 25343
        1033: data_ff <= 24'hFFC98A; // -13942
        1034: data_ff <= 24'h001BD3; // 7123
        1035: data_ff <= 24'hFFF30F; // -3313
        1036: data_ff <= 24'h000553; // 1363
        1037: data_ff <= 24'hFFFE2A; // -470
        1038: data_ff <= 24'h000076; // 118
        1039: data_ff <= 24'hFFFFF4; // -12
        1040: data_ff <= 24'h20E2F4; // 2155252
        1041: data_ff <= 24'hF458F2; // -763662
        1042: data_ff <= 24'h06862B; // 427563
        1043: data_ff <= 24'hFBE717; // -268521
        1044: data_ff <= 24'h02A88A; // 174218
        1045: data_ff <= 24'hFE4755; // -112811
        1046: data_ff <= 24'h011750; // 71504
        1047: data_ff <= 24'hFF5510; // -43760
        1048: data_ff <= 24'h0063CF; // 25551
        1049: data_ff <= 24'hFFC913; // -14061
        1050: data_ff <= 24'h001C12; // 7186
        1051: data_ff <= 24'hFFF2EF; // -3345
        1052: data_ff <= 24'h000561; // 1377
        1053: data_ff <= 24'hFFFE25; // -475
        1054: data_ff <= 24'h000078; // 120
        1055: data_ff <= 24'hFFFFF4; // -12
        1056: data_ff <= 24'h216CCA; // 2190538
        1057: data_ff <= 24'hF43BF6; // -771082
        1058: data_ff <= 24'h069410; // 431120
        1059: data_ff <= 24'hFBDEEC; // -270612
        1060: data_ff <= 24'h02ADB0; // 175536
        1061: data_ff <= 24'hFE4407; // -113657
        1062: data_ff <= 24'h01196A; // 72042
        1063: data_ff <= 24'hFF53C2; // -44094
        1064: data_ff <= 24'h006497; // 25751
        1065: data_ff <= 24'hFFC8A1; // -14175
        1066: data_ff <= 24'h001C4F; // 7247
        1067: data_ff <= 24'hFFF2D1; // -3375
        1068: data_ff <= 24'h00056E; // 1390
        1069: data_ff <= 24'hFFFE1F; // -481
        1070: data_ff <= 24'h00007A; // 122
        1071: data_ff <= 24'hFFFFF3; // -13
        1072: data_ff <= 24'h21F649; // 2225737
        1073: data_ff <= 24'hF41FE7; // -778265
        1074: data_ff <= 24'h06A163; // 434531
        1075: data_ff <= 24'hFBD71F; // -272609
        1076: data_ff <= 24'h02B298; // 176792
        1077: data_ff <= 24'hFE40E1; // -114463
        1078: data_ff <= 24'h011B6C; // 72556
        1079: data_ff <= 24'hFF5283; // -44413
        1080: data_ff <= 24'h006556; // 25942
        1081: data_ff <= 24'hFFC834; // -14284
        1082: data_ff <= 24'h001C89; // 7305
        1083: data_ff <= 24'hFFF2B4; // -3404
        1084: data_ff <= 24'h00057B; // 1403
        1085: data_ff <= 24'hFFFE1A; // -486
        1086: data_ff <= 24'h00007B; // 123
        1087: data_ff <= 24'hFFFFF3; // -13
        1088: data_ff <= 24'h227F69; // 2260841
        1089: data_ff <= 24'hF404C8; // -785208
        1090: data_ff <= 24'h06AE22; // 437794
        1091: data_ff <= 24'hFBCFB2; // -274510
        1092: data_ff <= 24'h02B742; // 177986
        1093: data_ff <= 24'hFE3DE4; // -115228
        1094: data_ff <= 24'h011D53; // 73043
        1095: data_ff <= 24'hFF5154; // -44716
        1096: data_ff <= 24'h00660D; // 26125
        1097: data_ff <= 24'hFFC7CC; // -14388
        1098: data_ff <= 24'h001CC1; // 7361
        1099: data_ff <= 24'hFFF299; // -3431
        1100: data_ff <= 24'h000588; // 1416
        1101: data_ff <= 24'hFFFE15; // -491
        1102: data_ff <= 24'h00007D; // 125
        1103: data_ff <= 24'hFFFFF3; // -13
        1104: data_ff <= 24'h230824; // 2295844
        1105: data_ff <= 24'hF3EA9E; // -791906
        1106: data_ff <= 24'h06BA4A; // 440906
        1107: data_ff <= 24'hFBC8A6; // -276314
        1108: data_ff <= 24'h02BBAC; // 179116
        1109: data_ff <= 24'hFE3B10; // -115952
        1110: data_ff <= 24'h011F21; // 73505
        1111: data_ff <= 24'hFF5034; // -45004
        1112: data_ff <= 24'h0066B9; // 26297
        1113: data_ff <= 24'hFFC769; // -14487
        1114: data_ff <= 24'h001CF7; // 7415
        1115: data_ff <= 24'hFFF27E; // -3458
        1116: data_ff <= 24'h000594; // 1428
        1117: data_ff <= 24'hFFFE10; // -496
        1118: data_ff <= 24'h00007E; // 126
        1119: data_ff <= 24'hFFFFF3; // -13
        1120: data_ff <= 24'h239070; // 2330736
        1121: data_ff <= 24'hF3D16E; // -798354
        1122: data_ff <= 24'h06C5D9; // 443865
        1123: data_ff <= 24'hFBC1FC; // -278020
        1124: data_ff <= 24'h02BFD7; // 180183
        1125: data_ff <= 24'hFE3865; // -116635
        1126: data_ff <= 24'h0120D4; // 73940
        1127: data_ff <= 24'hFF4F25; // -45275
        1128: data_ff <= 24'h00675D; // 26461
        1129: data_ff <= 24'hFFC70B; // -14581
        1130: data_ff <= 24'h001D29; // 7465
        1131: data_ff <= 24'hFFF264; // -3484
        1132: data_ff <= 24'h00059F; // 1439
        1133: data_ff <= 24'hFFFE0C; // -500
        1134: data_ff <= 24'h000080; // 128
        1135: data_ff <= 24'hFFFFF2; // -14
        1136: data_ff <= 24'h241847; // 2365511
        1137: data_ff <= 24'hF3B93D; // -804547
        1138: data_ff <= 24'h06D0CE; // 446670
        1139: data_ff <= 24'hFBBBB5; // -279627
        1140: data_ff <= 24'h02C3C0; // 181184
        1141: data_ff <= 24'hFE35E4; // -117276
        1142: data_ff <= 24'h01226D; // 74349
        1143: data_ff <= 24'hFF4E25; // -45531
        1144: data_ff <= 24'h0067F7; // 26615
        1145: data_ff <= 24'hFFC6B2; // -14670
        1146: data_ff <= 24'h001D5A; // 7514
        1147: data_ff <= 24'hFFF24C; // -3508
        1148: data_ff <= 24'h0005AB; // 1451
        1149: data_ff <= 24'hFFFE07; // -505
        1150: data_ff <= 24'h000081; // 129
        1151: data_ff <= 24'hFFFFF2; // -14
        1152: data_ff <= 24'h249FA1; // 2400161
        1153: data_ff <= 24'hF3A20F; // -810481
        1154: data_ff <= 24'h06DB26; // 449318
        1155: data_ff <= 24'hFBB5D2; // -281134
        1156: data_ff <= 24'h02C767; // 182119
        1157: data_ff <= 24'hFE338E; // -117874
        1158: data_ff <= 24'h0123EA; // 74730
        1159: data_ff <= 24'hFF4D36; // -45770
        1160: data_ff <= 24'h006888; // 26760
        1161: data_ff <= 24'hFFC65F; // -14753
        1162: data_ff <= 24'h001D87; // 7559
        1163: data_ff <= 24'hFFF235; // -3531
        1164: data_ff <= 24'h0005B5; // 1461
        1165: data_ff <= 24'hFFFE03; // -509
        1166: data_ff <= 24'h000083; // 131
        1167: data_ff <= 24'hFFFFF2; // -14
        1168: data_ff <= 24'h252676; // 2434678
        1169: data_ff <= 24'hF38BE8; // -816152
        1170: data_ff <= 24'h06E4DF; // 451807
        1171: data_ff <= 24'hFBB056; // -282538
        1172: data_ff <= 24'h02CACD; // 182989
        1173: data_ff <= 24'hFE3163; // -118429
        1174: data_ff <= 24'h01254D; // 75085
        1175: data_ff <= 24'hFF4C58; // -45992
        1176: data_ff <= 24'h00690F; // 26895
        1177: data_ff <= 24'hFFC610; // -14832
        1178: data_ff <= 24'h001DB2; // 7602
        1179: data_ff <= 24'hFFF21F; // -3553
        1180: data_ff <= 24'h0005BF; // 1471
        1181: data_ff <= 24'hFFFDFF; // -513
        1182: data_ff <= 24'h000084; // 132
        1183: data_ff <= 24'hFFFFF1; // -15
        1184: data_ff <= 24'h25ACBF; // 2469055
        1185: data_ff <= 24'hF376CE; // -821554
        1186: data_ff <= 24'h06EDF8; // 454136
        1187: data_ff <= 24'hFBAB40; // -283840
        1188: data_ff <= 24'h02CDEF; // 183791
        1189: data_ff <= 24'hFE2F64; // -118940
        1190: data_ff <= 24'h012694; // 75412
        1191: data_ff <= 24'hFF4B8B; // -46197
        1192: data_ff <= 24'h00698C; // 27020
        1193: data_ff <= 24'hFFC5C7; // -14905
        1194: data_ff <= 24'h001DDB; // 7643
        1195: data_ff <= 24'hFFF20A; // -3574
        1196: data_ff <= 24'h0005C9; // 1481
        1197: data_ff <= 24'hFFFDFB; // -517
        1198: data_ff <= 24'h000086; // 134
        1199: data_ff <= 24'hFFFFF1; // -15
        1200: data_ff <= 24'h263274; // 2503284
        1201: data_ff <= 24'hF362C4; // -826684
        1202: data_ff <= 24'h06F66E; // 456302
        1203: data_ff <= 24'hFBA691; // -285039
        1204: data_ff <= 24'h02D0CE; // 184526
        1205: data_ff <= 24'hFE2D91; // -119407
        1206: data_ff <= 24'h0127BF; // 75711
        1207: data_ff <= 24'hFF4ACE; // -46386
        1208: data_ff <= 24'h0069FF; // 27135
        1209: data_ff <= 24'hFFC584; // -14972
        1210: data_ff <= 24'h001E00; // 7680
        1211: data_ff <= 24'hFFF1F7; // -3593
        1212: data_ff <= 24'h0005D2; // 1490
        1213: data_ff <= 24'hFFFDF7; // -521
        1214: data_ff <= 24'h000087; // 135
        1215: data_ff <= 24'hFFFFF1; // -15
        1216: data_ff <= 24'h26B78E; // 2537358
        1217: data_ff <= 24'hF34FCE; // -831538
        1218: data_ff <= 24'h06FE3F; // 458303
        1219: data_ff <= 24'hFBA24C; // -286132
        1220: data_ff <= 24'h02D368; // 185192
        1221: data_ff <= 24'hFE2BE9; // -119831
        1222: data_ff <= 24'h0128CD; // 75981
        1223: data_ff <= 24'hFF4A23; // -46557
        1224: data_ff <= 24'h006A68; // 27240
        1225: data_ff <= 24'hFFC546; // -15034
        1226: data_ff <= 24'h001E23; // 7715
        1227: data_ff <= 24'hFFF1E5; // -3611
        1228: data_ff <= 24'h0005DB; // 1499
        1229: data_ff <= 24'hFFFDF3; // -525
        1230: data_ff <= 24'h000088; // 136
        1231: data_ff <= 24'hFFFFF1; // -15
        1232: data_ff <= 24'h273C04; // 2571268
        1233: data_ff <= 24'hF33DF1; // -836111
        1234: data_ff <= 24'h07056A; // 460138
        1235: data_ff <= 24'hFB9E70; // -287120
        1236: data_ff <= 24'h02D5BD; // 185789
        1237: data_ff <= 24'hFE2A6F; // -120209
        1238: data_ff <= 24'h0129C0; // 76224
        1239: data_ff <= 24'hFF4989; // -46711
        1240: data_ff <= 24'h006AC7; // 27335
        1241: data_ff <= 24'hFFC50D; // -15091
        1242: data_ff <= 24'h001E43; // 7747
        1243: data_ff <= 24'hFFF1D4; // -3628
        1244: data_ff <= 24'h0005E3; // 1507
        1245: data_ff <= 24'hFFFDF0; // -528
        1246: data_ff <= 24'h00008A; // 138
        1247: data_ff <= 24'hFFFFF0; // -16
        1248: data_ff <= 24'h27BFD0; // 2605008
        1249: data_ff <= 24'hF32D32; // -840398
        1250: data_ff <= 24'h070BED; // 461805
        1251: data_ff <= 24'hFB9B00; // -288000
        1252: data_ff <= 24'h02D7CC; // 186316
        1253: data_ff <= 24'hFE2922; // -120542
        1254: data_ff <= 24'h012A96; // 76438
        1255: data_ff <= 24'hFF4901; // -46847
        1256: data_ff <= 24'h006B1C; // 27420
        1257: data_ff <= 24'hFFC4DA; // -15142
        1258: data_ff <= 24'h001E60; // 7776
        1259: data_ff <= 24'hFFF1C5; // -3643
        1260: data_ff <= 24'h0005EA; // 1514
        1261: data_ff <= 24'hFFFDED; // -531
        1262: data_ff <= 24'h00008B; // 139
        1263: data_ff <= 24'hFFFFF0; // -16
        1264: data_ff <= 24'h2842EA; // 2638570
        1265: data_ff <= 24'hF31D94; // -844396
        1266: data_ff <= 24'h0711C7; // 463303
        1267: data_ff <= 24'hFB97FB; // -288773
        1268: data_ff <= 24'h02D995; // 186773
        1269: data_ff <= 24'hFE2802; // -120830
        1270: data_ff <= 24'h012B4F; // 76623
        1271: data_ff <= 24'hFF488B; // -46965
        1272: data_ff <= 24'h006B67; // 27495
        1273: data_ff <= 24'hFFC4AD; // -15187
        1274: data_ff <= 24'h001E7A; // 7802
        1275: data_ff <= 24'hFFF1B7; // -3657
        1276: data_ff <= 24'h0005F1; // 1521
        1277: data_ff <= 24'hFFFDEA; // -534
        1278: data_ff <= 24'h00008C; // 140
        1279: data_ff <= 24'hFFFFF0; // -16
        1280: data_ff <= 24'h28C54B; // 2671947
        1281: data_ff <= 24'hF30F1B; // -848101
        1282: data_ff <= 24'h0716F4; // 464628
        1283: data_ff <= 24'hFB9563; // -289437
        1284: data_ff <= 24'h02DB18; // 187160
        1285: data_ff <= 24'hFE2711; // -121071
        1286: data_ff <= 24'h012BEA; // 76778
        1287: data_ff <= 24'hFF4826; // -47066
        1288: data_ff <= 24'h006BA7; // 27559
        1289: data_ff <= 24'hFFC486; // -15226
        1290: data_ff <= 24'h001E91; // 7825
        1291: data_ff <= 24'hFFF1AA; // -3670
        1292: data_ff <= 24'h0005F8; // 1528
        1293: data_ff <= 24'hFFFDE7; // -537
        1294: data_ff <= 24'h00008D; // 141
        1295: data_ff <= 24'hFFFFEF; // -17
        1296: data_ff <= 24'h2946EA; // 2705130
        1297: data_ff <= 24'hF301CB; // -851509
        1298: data_ff <= 24'h071B75; // 465781
        1299: data_ff <= 24'hFB9338; // -289992
        1300: data_ff <= 24'h02DC53; // 187475
        1301: data_ff <= 24'hFE264D; // -121267
        1302: data_ff <= 24'h012C69; // 76905
        1303: data_ff <= 24'hFF47D3; // -47149
        1304: data_ff <= 24'h006BDC; // 27612
        1305: data_ff <= 24'hFFC464; // -15260
        1306: data_ff <= 24'h001EA5; // 7845
        1307: data_ff <= 24'hFFF19F; // -3681
        1308: data_ff <= 24'h0005FD; // 1533
        1309: data_ff <= 24'hFFFDE4; // -540
        1310: data_ff <= 24'h00008E; // 142
        1311: data_ff <= 24'hFFFFEF; // -17
        1312: data_ff <= 24'h29C7C1; // 2738113
        1313: data_ff <= 24'hF2F5A9; // -854615
        1314: data_ff <= 24'h071F47; // 466759
        1315: data_ff <= 24'hFB917C; // -290436
        1316: data_ff <= 24'h02DD46; // 187718
        1317: data_ff <= 24'hFE25B8; // -121416
        1318: data_ff <= 24'h012CC9; // 77001
        1319: data_ff <= 24'hFF4793; // -47213
        1320: data_ff <= 24'h006C07; // 27655
        1321: data_ff <= 24'hFFC449; // -15287
        1322: data_ff <= 24'h001EB6; // 7862
        1323: data_ff <= 24'hFFF195; // -3691
        1324: data_ff <= 24'h000603; // 1539
        1325: data_ff <= 24'hFFFDE2; // -542
        1326: data_ff <= 24'h00008F; // 143
        1327: data_ff <= 24'hFFFFEF; // -17
        1328: data_ff <= 24'h2A47C8; // 2770888
        1329: data_ff <= 24'hF2EAB9; // -857415
        1330: data_ff <= 24'h072269; // 467561
        1331: data_ff <= 24'hFB902F; // -290769
        1332: data_ff <= 24'h02DDF1; // 187889
        1333: data_ff <= 24'hFE2553; // -121517
        1334: data_ff <= 24'h012D0C; // 77068
        1335: data_ff <= 24'hFF4765; // -47259
        1336: data_ff <= 24'h006C27; // 27687
        1337: data_ff <= 24'hFFC433; // -15309
        1338: data_ff <= 24'h001EC4; // 7876
        1339: data_ff <= 24'hFFF18D; // -3699
        1340: data_ff <= 24'h000607; // 1543
        1341: data_ff <= 24'hFFFDDF; // -545
        1342: data_ff <= 24'h000090; // 144
        1343: data_ff <= 24'hFFFFEF; // -17
        1344: data_ff <= 24'h2AC6F8; // 2803448
        1345: data_ff <= 24'hF2E0FD; // -859907
        1346: data_ff <= 24'h0724D9; // 468185
        1347: data_ff <= 24'hFB8F51; // -290991
        1348: data_ff <= 24'h02DE54; // 187988
        1349: data_ff <= 24'hFE251C; // -121572
        1350: data_ff <= 24'h012D31; // 77105
        1351: data_ff <= 24'hFF4749; // -47287
        1352: data_ff <= 24'h006C3C; // 27708
        1353: data_ff <= 24'hFFC423; // -15325
        1354: data_ff <= 24'h001ECF; // 7887
        1355: data_ff <= 24'hFFF186; // -3706
        1356: data_ff <= 24'h00060B; // 1547
        1357: data_ff <= 24'hFFFDDD; // -547
        1358: data_ff <= 24'h000091; // 145
        1359: data_ff <= 24'hFFFFEE; // -18
        1360: data_ff <= 24'h2B4549; // 2835785
        1361: data_ff <= 24'hF2D87A; // -862086
        1362: data_ff <= 24'h072697; // 468631
        1363: data_ff <= 24'hFB8EE5; // -291099
        1364: data_ff <= 24'h02DE6D; // 188013
        1365: data_ff <= 24'hFE2515; // -121579
        1366: data_ff <= 24'h012D37; // 77111
        1367: data_ff <= 24'hFF4740; // -47296
        1368: data_ff <= 24'h006C46; // 27718
        1369: data_ff <= 24'hFFC41A; // -15334
        1370: data_ff <= 24'h001ED6; // 7894
        1371: data_ff <= 24'hFFF180; // -3712
        1372: data_ff <= 24'h00060F; // 1551
        1373: data_ff <= 24'hFFFDDC; // -548
        1374: data_ff <= 24'h000092; // 146
        1375: data_ff <= 24'hFFFFEE; // -18
        1376: data_ff <= 24'h2BC2B5; // 2867893
        1377: data_ff <= 24'hF2D134; // -863948
        1378: data_ff <= 24'h0727A0; // 468896
        1379: data_ff <= 24'hFB8EEA; // -291094
        1380: data_ff <= 24'h02DE3D; // 187965
        1381: data_ff <= 24'hFE253E; // -121538
        1382: data_ff <= 24'h012D20; // 77088
        1383: data_ff <= 24'hFF474A; // -47286
        1384: data_ff <= 24'h006C45; // 27717
        1385: data_ff <= 24'hFFC416; // -15338
        1386: data_ff <= 24'h001EDB; // 7899
        1387: data_ff <= 24'hFFF17C; // -3716
        1388: data_ff <= 24'h000611; // 1553
        1389: data_ff <= 24'hFFFDDA; // -550
        1390: data_ff <= 24'h000093; // 147
        1391: data_ff <= 24'hFFFFEE; // -18
        1392: data_ff <= 24'h2C3F34; // 2899764
        1393: data_ff <= 24'hF2CB2F; // -865489
        1394: data_ff <= 24'h0727F3; // 468979
        1395: data_ff <= 24'hFB8F60; // -290976
        1396: data_ff <= 24'h02DDC2; // 187842
        1397: data_ff <= 24'hFE2596; // -121450
        1398: data_ff <= 24'h012CE9; // 77033
        1399: data_ff <= 24'hFF4767; // -47257
        1400: data_ff <= 24'h006C39; // 27705
        1401: data_ff <= 24'hFFC419; // -15335
        1402: data_ff <= 24'h001EDD; // 7901
        1403: data_ff <= 24'hFFF17A; // -3718
        1404: data_ff <= 24'h000614; // 1556
        1405: data_ff <= 24'hFFFDD9; // -551
        1406: data_ff <= 24'h000093; // 147
        1407: data_ff <= 24'hFFFFEE; // -18
        1408: data_ff <= 24'h2CBABE; // 2931390
        1409: data_ff <= 24'hF2C66D; // -866707
        1410: data_ff <= 24'h072790; // 468880
        1411: data_ff <= 24'hFB9049; // -290743
        1412: data_ff <= 24'h02DCFD; // 187645
        1413: data_ff <= 24'hFE261F; // -121313
        1414: data_ff <= 24'h012C94; // 76948
        1415: data_ff <= 24'hFF4796; // -47210
        1416: data_ff <= 24'h006C22; // 27682
        1417: data_ff <= 24'hFFC422; // -15326
        1418: data_ff <= 24'h001EDB; // 7899
        1419: data_ff <= 24'hFFF179; // -3719
        1420: data_ff <= 24'h000615; // 1557
        1421: data_ff <= 24'hFFFDD7; // -553
        1422: data_ff <= 24'h000094; // 148
        1423: data_ff <= 24'hFFFFED; // -19
        1424: data_ff <= 24'h2D354D; // 2962765
        1425: data_ff <= 24'hF2C2F2; // -867598
        1426: data_ff <= 24'h072675; // 468597
        1427: data_ff <= 24'hFB91A6; // -290394
        1428: data_ff <= 24'h02DBEE; // 187374
        1429: data_ff <= 24'hFE26D9; // -121127
        1430: data_ff <= 24'h012C20; // 76832
        1431: data_ff <= 24'hFF47D9; // -47143
        1432: data_ff <= 24'h006C00; // 27648
        1433: data_ff <= 24'hFFC431; // -15311
        1434: data_ff <= 24'h001ED6; // 7894
        1435: data_ff <= 24'hFFF179; // -3719
        1436: data_ff <= 24'h000616; // 1558
        1437: data_ff <= 24'hFFFDD7; // -553
        1438: data_ff <= 24'h000094; // 148
        1439: data_ff <= 24'hFFFFED; // -19
        1440: data_ff <= 24'h2DAEDA; // 2993882
        1441: data_ff <= 24'hF2C0C3; // -868157
        1442: data_ff <= 24'h0724A1; // 468129
        1443: data_ff <= 24'hFB9375; // -289931
        1444: data_ff <= 24'h02DA94; // 187028
        1445: data_ff <= 24'hFE27C3; // -120893
        1446: data_ff <= 24'h012B8D; // 76685
        1447: data_ff <= 24'hFF482E; // -47058
        1448: data_ff <= 24'h006BD3; // 27603
        1449: data_ff <= 24'hFFC446; // -15290
        1450: data_ff <= 24'h001ECD; // 7885
        1451: data_ff <= 24'hFFF17B; // -3717
        1452: data_ff <= 24'h000616; // 1558
        1453: data_ff <= 24'hFFFDD6; // -554
        1454: data_ff <= 24'h000095; // 149
        1455: data_ff <= 24'hFFFFED; // -19
        1456: data_ff <= 24'h2E275D; // 3024733
        1457: data_ff <= 24'hF2BFE1; // -868383
        1458: data_ff <= 24'h072213; // 467475
        1459: data_ff <= 24'hFB95B9; // -289351
        1460: data_ff <= 24'h02D8EE; // 186606
        1461: data_ff <= 24'hFE28DD; // -120611
        1462: data_ff <= 24'h012ADB; // 76507
        1463: data_ff <= 24'hFF4897; // -46953
        1464: data_ff <= 24'h006B9A; // 27546
        1465: data_ff <= 24'hFFC462; // -15262
        1466: data_ff <= 24'h001EC2; // 7874
        1467: data_ff <= 24'hFFF17F; // -3713
        1468: data_ff <= 24'h000616; // 1558
        1469: data_ff <= 24'hFFFDD5; // -555
        1470: data_ff <= 24'h000095; // 149
        1471: data_ff <= 24'hFFFFED; // -19
        1472: data_ff <= 24'h2E9ECF; // 3055311
        1473: data_ff <= 24'hF2C051; // -868271
        1474: data_ff <= 24'h071ECA; // 466634
        1475: data_ff <= 24'hFB9872; // -288654
        1476: data_ff <= 24'h02D6FD; // 186109
        1477: data_ff <= 24'hFE2A29; // -120279
        1478: data_ff <= 24'h012A09; // 76297
        1479: data_ff <= 24'hFF4913; // -46829
        1480: data_ff <= 24'h006B55; // 27477
        1481: data_ff <= 24'hFFC484; // -15228
        1482: data_ff <= 24'h001EB3; // 7859
        1483: data_ff <= 24'hFFF184; // -3708
        1484: data_ff <= 24'h000615; // 1557
        1485: data_ff <= 24'hFFFDD5; // -555
        1486: data_ff <= 24'h000096; // 150
        1487: data_ff <= 24'hFFFFED; // -19
        1488: data_ff <= 24'h2F152A; // 3085610
        1489: data_ff <= 24'hF2C215; // -867819
        1490: data_ff <= 24'h071AC5; // 465605
        1491: data_ff <= 24'hFB9B9F; // -287841
        1492: data_ff <= 24'h02D4C1; // 185537
        1493: data_ff <= 24'hFE2BA6; // -119898
        1494: data_ff <= 24'h012919; // 76057
        1495: data_ff <= 24'hFF49A3; // -46685
        1496: data_ff <= 24'h006B06; // 27398
        1497: data_ff <= 24'hFFC4AD; // -15187
        1498: data_ff <= 24'h001EA1; // 7841
        1499: data_ff <= 24'hFFF18B; // -3701
        1500: data_ff <= 24'h000613; // 1555
        1501: data_ff <= 24'hFFFDD5; // -555
        1502: data_ff <= 24'h000096; // 150
        1503: data_ff <= 24'hFFFFEC; // -20
        1504: data_ff <= 24'h2F8A66; // 3115622
        1505: data_ff <= 24'hF2C532; // -867022
        1506: data_ff <= 24'h071603; // 464387
        1507: data_ff <= 24'hFB9F41; // -286911
        1508: data_ff <= 24'h02D238; // 184888
        1509: data_ff <= 24'hFE2D55; // -119467
        1510: data_ff <= 24'h012808; // 75784
        1511: data_ff <= 24'hFF4A46; // -46522
        1512: data_ff <= 24'h006AAA; // 27306
        1513: data_ff <= 24'hFFC4DC; // -15140
        1514: data_ff <= 24'h001E8B; // 7819
        1515: data_ff <= 24'hFFF193; // -3693
        1516: data_ff <= 24'h000610; // 1552
        1517: data_ff <= 24'hFFFDD6; // -554
        1518: data_ff <= 24'h000096; // 150
        1519: data_ff <= 24'hFFFFEC; // -20
        1520: data_ff <= 24'h2FFE7D; // 3145341
        1521: data_ff <= 24'hF2C9A9; // -865879
        1522: data_ff <= 24'h071084; // 462980
        1523: data_ff <= 24'hFBA359; // -285863
        1524: data_ff <= 24'h02CF64; // 184164
        1525: data_ff <= 24'hFE2F34; // -118988
        1526: data_ff <= 24'h0126D9; // 75481
        1527: data_ff <= 24'hFF4AFC; // -46340
        1528: data_ff <= 24'h006A44; // 27204
        1529: data_ff <= 24'hFFC511; // -15087
        1530: data_ff <= 24'h001E72; // 7794
        1531: data_ff <= 24'hFFF19E; // -3682
        1532: data_ff <= 24'h00060D; // 1549
        1533: data_ff <= 24'hFFFDD6; // -554
        1534: data_ff <= 24'h000097; // 151
        1535: data_ff <= 24'hFFFFEC; // -20
        1536: data_ff <= 24'h307168; // 3174760
        1537: data_ff <= 24'hF2CF7E; // -864386
        1538: data_ff <= 24'h070A46; // 461382
        1539: data_ff <= 24'hFBA7E7; // -284697
        1540: data_ff <= 24'h02CC44; // 183364
        1541: data_ff <= 24'hFE3145; // -118459
        1542: data_ff <= 24'h012589; // 75145
        1543: data_ff <= 24'hFF4BC6; // -46138
        1544: data_ff <= 24'h0069D1; // 27089
        1545: data_ff <= 24'hFFC54D; // -15027
        1546: data_ff <= 24'h001E56; // 7766
        1547: data_ff <= 24'hFFF1A9; // -3671
        1548: data_ff <= 24'h000609; // 1545
        1549: data_ff <= 24'hFFFDD7; // -553
        1550: data_ff <= 24'h000097; // 151
        1551: data_ff <= 24'hFFFFEC; // -20
        1552: data_ff <= 24'h30E321; // 3203873
        1553: data_ff <= 24'hF2D6B3; // -862541
        1554: data_ff <= 24'h07034A; // 459594
        1555: data_ff <= 24'hFBACEA; // -283414
        1556: data_ff <= 24'h02C8D7; // 182487
        1557: data_ff <= 24'hFE3388; // -117880
        1558: data_ff <= 24'h01241B; // 74779
        1559: data_ff <= 24'hFF4CA4; // -45916
        1560: data_ff <= 24'h006953; // 26963
        1561: data_ff <= 24'hFFC58F; // -14961
        1562: data_ff <= 24'h001E36; // 7734
        1563: data_ff <= 24'hFFF1B7; // -3657
        1564: data_ff <= 24'h000605; // 1541
        1565: data_ff <= 24'hFFFDD8; // -552
        1566: data_ff <= 24'h000097; // 151
        1567: data_ff <= 24'hFFFFEC; // -20
        1568: data_ff <= 24'h31539F; // 3232671
        1569: data_ff <= 24'hF2DF4C; // -860340
        1570: data_ff <= 24'h06FB8E; // 457614
        1571: data_ff <= 24'hFBB264; // -282012
        1572: data_ff <= 24'h02C51E; // 181534
        1573: data_ff <= 24'hFE35FC; // -117252
        1574: data_ff <= 24'h01228C; // 74380
        1575: data_ff <= 24'hFF4D95; // -45675
        1576: data_ff <= 24'h0068C9; // 26825
        1577: data_ff <= 24'hFFC5D8; // -14888
        1578: data_ff <= 24'h001E13; // 7699
        1579: data_ff <= 24'hFFF1C6; // -3642
        1580: data_ff <= 24'h0005FF; // 1535
        1581: data_ff <= 24'hFFFDD9; // -551
        1582: data_ff <= 24'h000097; // 151
        1583: data_ff <= 24'hFFFFEB; // -21
        1584: data_ff <= 24'h31C2DE; // 3261150
        1585: data_ff <= 24'hF2E94B; // -857781
        1586: data_ff <= 24'h06F313; // 455443
        1587: data_ff <= 24'hFBB854; // -280492
        1588: data_ff <= 24'h02C119; // 180505
        1589: data_ff <= 24'hFE38A1; // -116575
        1590: data_ff <= 24'h0120DE; // 73950
        1591: data_ff <= 24'hFF4E9A; // -45414
        1592: data_ff <= 24'h006834; // 26676
        1593: data_ff <= 24'hFFC628; // -14808
        1594: data_ff <= 24'h001DEC; // 7660
        1595: data_ff <= 24'hFFF1D6; // -3626
        1596: data_ff <= 24'h0005F9; // 1529
        1597: data_ff <= 24'hFFFDDB; // -549
        1598: data_ff <= 24'h000097; // 151
        1599: data_ff <= 24'hFFFFEB; // -21
        1600: data_ff <= 24'h3230D6; // 3289302
        1601: data_ff <= 24'hF2F4B3; // -854861
        1602: data_ff <= 24'h06E9D6; // 453078
        1603: data_ff <= 24'hFBBEBA; // -278854
        1604: data_ff <= 24'h02BCC7; // 179399
        1605: data_ff <= 24'hFE3B79; // -115847
        1606: data_ff <= 24'h011F10; // 73488
        1607: data_ff <= 24'hFF4FB3; // -45133
        1608: data_ff <= 24'h006793; // 26515
        1609: data_ff <= 24'hFFC67E; // -14722
        1610: data_ff <= 24'h001DC2; // 7618
        1611: data_ff <= 24'hFFF1E9; // -3607
        1612: data_ff <= 24'h0005F3; // 1523
        1613: data_ff <= 24'hFFFDDD; // -547
        1614: data_ff <= 24'h000097; // 151
        1615: data_ff <= 24'hFFFFEB; // -21
        1616: data_ff <= 24'h329D81; // 3317121
        1617: data_ff <= 24'hF30186; // -851578
        1618: data_ff <= 24'h06DFDA; // 450522
        1619: data_ff <= 24'hFBC596; // -277098
        1620: data_ff <= 24'h02B829; // 178217
        1621: data_ff <= 24'hFE3E81; // -115071
        1622: data_ff <= 24'h011D22; // 72994
        1623: data_ff <= 24'hFF50DF; // -44833
        1624: data_ff <= 24'h0066E6; // 26342
        1625: data_ff <= 24'hFFC6DB; // -14629
        1626: data_ff <= 24'h001D94; // 7572
        1627: data_ff <= 24'hFFF1FD; // -3587
        1628: data_ff <= 24'h0005EB; // 1515
        1629: data_ff <= 24'hFFFDDF; // -545
        1630: data_ff <= 24'h000096; // 150
        1631: data_ff <= 24'hFFFFEB; // -21
        1632: data_ff <= 24'h3308D8; // 3344600
        1633: data_ff <= 24'hF30FC8; // -847928
        1634: data_ff <= 24'h06D51C; // 447772
        1635: data_ff <= 24'hFBCCE9; // -275223
        1636: data_ff <= 24'h02B33F; // 176959
        1637: data_ff <= 24'hFE41BC; // -114244
        1638: data_ff <= 24'h011B15; // 72469
        1639: data_ff <= 24'hFF521F; // -44513
        1640: data_ff <= 24'h00662E; // 26158
        1641: data_ff <= 24'hFFC73E; // -14530
        1642: data_ff <= 24'h001D63; // 7523
        1643: data_ff <= 24'hFFF212; // -3566
        1644: data_ff <= 24'h0005E3; // 1507
        1645: data_ff <= 24'hFFFDE1; // -543
        1646: data_ff <= 24'h000096; // 150
        1647: data_ff <= 24'hFFFFEB; // -21
        1648: data_ff <= 24'h3372D6; // 3371734
        1649: data_ff <= 24'hF31F79; // -843911
        1650: data_ff <= 24'h06C99D; // 444829
        1651: data_ff <= 24'hFBD4B3; // -273229
        1652: data_ff <= 24'h02AE09; // 175625
        1653: data_ff <= 24'hFE4527; // -113369
        1654: data_ff <= 24'h0118E8; // 71912
        1655: data_ff <= 24'hFF5372; // -44174
        1656: data_ff <= 24'h00656A; // 25962
        1657: data_ff <= 24'hFFC7A8; // -14424
        1658: data_ff <= 24'h001D2F; // 7471
        1659: data_ff <= 24'hFFF22A; // -3542
        1660: data_ff <= 24'h0005DA; // 1498
        1661: data_ff <= 24'hFFFDE4; // -540
        1662: data_ff <= 24'h000095; // 149
        1663: data_ff <= 24'hFFFFEB; // -21
        1664: data_ff <= 24'h33DB73; // 3398515
        1665: data_ff <= 24'hF3309D; // -839523
        1666: data_ff <= 24'h06BD5C; // 441692
        1667: data_ff <= 24'hFBDCF2; // -271118
        1668: data_ff <= 24'h02A886; // 174214
        1669: data_ff <= 24'hFE48C4; // -112444
        1670: data_ff <= 24'h01169B; // 71323
        1671: data_ff <= 24'hFF54D9; // -43815
        1672: data_ff <= 24'h00649A; // 25754
        1673: data_ff <= 24'hFFC819; // -14311
        1674: data_ff <= 24'h001CF6; // 7414
        1675: data_ff <= 24'hFFF243; // -3517
        1676: data_ff <= 24'h0005D0; // 1488
        1677: data_ff <= 24'hFFFDE7; // -537
        1678: data_ff <= 24'h000095; // 149
        1679: data_ff <= 24'hFFFFEB; // -21
        1680: data_ff <= 24'h3442AA; // 3424938
        1681: data_ff <= 24'hF34335; // -834763
        1682: data_ff <= 24'h06B05A; // 438362
        1683: data_ff <= 24'hFBE5A7; // -268889
        1684: data_ff <= 24'h02A2B8; // 172728
        1685: data_ff <= 24'hFE4C93; // -111469
        1686: data_ff <= 24'h01142F; // 70703
        1687: data_ff <= 24'hFF5654; // -43436
        1688: data_ff <= 24'h0063BE; // 25534
        1689: data_ff <= 24'hFFC890; // -14192
        1690: data_ff <= 24'h001CBB; // 7355
        1691: data_ff <= 24'hFFF25E; // -3490
        1692: data_ff <= 24'h0005C6; // 1478
        1693: data_ff <= 24'hFFFDEA; // -534
        1694: data_ff <= 24'h000094; // 148
        1695: data_ff <= 24'hFFFFEB; // -21
        1696: data_ff <= 24'h34A875; // 3450997
        1697: data_ff <= 24'hF35744; // -829628
        1698: data_ff <= 24'h06A296; // 434838
        1699: data_ff <= 24'hFBEED2; // -266542
        1700: data_ff <= 24'h029C9E; // 171166
        1701: data_ff <= 24'hFE5092; // -110446
        1702: data_ff <= 24'h0111A3; // 70051
        1703: data_ff <= 24'hFF57E3; // -43037
        1704: data_ff <= 24'h0062D7; // 25303
        1705: data_ff <= 24'hFFC90E; // -14066
        1706: data_ff <= 24'h001C7C; // 7292
        1707: data_ff <= 24'hFFF27A; // -3462
        1708: data_ff <= 24'h0005BB; // 1467
        1709: data_ff <= 24'hFFFDEE; // -530
        1710: data_ff <= 24'h000094; // 148
        1711: data_ff <= 24'hFFFFEB; // -21
        1712: data_ff <= 24'h350CCE; // 3476686
        1713: data_ff <= 24'hF36CCC; // -824116
        1714: data_ff <= 24'h069411; // 431121
        1715: data_ff <= 24'hFBF873; // -264077
        1716: data_ff <= 24'h029638; // 169528
        1717: data_ff <= 24'hFE54C3; // -109373
        1718: data_ff <= 24'h010EF8; // 69368
        1719: data_ff <= 24'hFF5985; // -42619
        1720: data_ff <= 24'h0061E4; // 25060
        1721: data_ff <= 24'hFFC992; // -13934
        1722: data_ff <= 24'h001C39; // 7225
        1723: data_ff <= 24'hFFF298; // -3432
        1724: data_ff <= 24'h0005AF; // 1455
        1725: data_ff <= 24'hFFFDF1; // -527
        1726: data_ff <= 24'h000093; // 147
        1727: data_ff <= 24'hFFFFEB; // -21
        1728: data_ff <= 24'h356FAD; // 3501997
        1729: data_ff <= 24'hF383CE; // -818226
        1730: data_ff <= 24'h0684CA; // 427210
        1731: data_ff <= 24'hFC0289; // -261495
        1732: data_ff <= 24'h028F87; // 167815
        1733: data_ff <= 24'hFE5925; // -108251
        1734: data_ff <= 24'h010C2E; // 68654
        1735: data_ff <= 24'hFF5B3A; // -42182
        1736: data_ff <= 24'h0060E5; // 24805
        1737: data_ff <= 24'hFFCA1E; // -13794
        1738: data_ff <= 24'h001BF3; // 7155
        1739: data_ff <= 24'hFFF2B8; // -3400
        1740: data_ff <= 24'h0005A2; // 1442
        1741: data_ff <= 24'hFFFDF5; // -523
        1742: data_ff <= 24'h000092; // 146
        1743: data_ff <= 24'hFFFFEB; // -21
        1744: data_ff <= 24'h35D10F; // 3526927
        1745: data_ff <= 24'hF39C4D; // -811955
        1746: data_ff <= 24'h0674C2; // 423106
        1747: data_ff <= 24'hFC0D14; // -258796
        1748: data_ff <= 24'h02888B; // 166027
        1749: data_ff <= 24'hFE5DB7; // -107081
        1750: data_ff <= 24'h010944; // 67908
        1751: data_ff <= 24'hFF5D04; // -41724
        1752: data_ff <= 24'h005FDB; // 24539
        1753: data_ff <= 24'hFFCAAF; // -13649
        1754: data_ff <= 24'h001BA9; // 7081
        1755: data_ff <= 24'hFFF2DA; // -3366
        1756: data_ff <= 24'h000595; // 1429
        1757: data_ff <= 24'hFFFDFA; // -518
        1758: data_ff <= 24'h000091; // 145
        1759: data_ff <= 24'hFFFFEB; // -21
        1760: data_ff <= 24'h3630ED; // 3551469
        1761: data_ff <= 24'hF3B64A; // -805302
        1762: data_ff <= 24'h0663F9; // 418809
        1763: data_ff <= 24'hFC1814; // -255980
        1764: data_ff <= 24'h028145; // 164165
        1765: data_ff <= 24'hFE627A; // -105862
        1766: data_ff <= 24'h01063B; // 67131
        1767: data_ff <= 24'hFF5EE0; // -41248
        1768: data_ff <= 24'h005EC5; // 24261
        1769: data_ff <= 24'hFFCB48; // -13496
        1770: data_ff <= 24'h001B5C; // 7004
        1771: data_ff <= 24'hFFF2FD; // -3331
        1772: data_ff <= 24'h000586; // 1414
        1773: data_ff <= 24'hFFFDFE; // -514
        1774: data_ff <= 24'h000090; // 144
        1775: data_ff <= 24'hFFFFEB; // -21
        1776: data_ff <= 24'h368F41; // 3575617
        1777: data_ff <= 24'hF3D1C7; // -798265
        1778: data_ff <= 24'h06526F; // 414319
        1779: data_ff <= 24'hFC2387; // -253049
        1780: data_ff <= 24'h0279B4; // 162228
        1781: data_ff <= 24'hFE676D; // -104595
        1782: data_ff <= 24'h010313; // 66323
        1783: data_ff <= 24'hFF60D0; // -40752
        1784: data_ff <= 24'h005DA3; // 23971
        1785: data_ff <= 24'hFFCBE7; // -13337
        1786: data_ff <= 24'h001B0B; // 6923
        1787: data_ff <= 24'hFFF323; // -3293
        1788: data_ff <= 24'h000577; // 1399
        1789: data_ff <= 24'hFFFE03; // -509
        1790: data_ff <= 24'h00008F; // 143
        1791: data_ff <= 24'hFFFFEB; // -21
        1792: data_ff <= 24'h36EC05; // 3599365
        1793: data_ff <= 24'hF3EEC5; // -790843
        1794: data_ff <= 24'h064026; // 409638
        1795: data_ff <= 24'hFC2F6F; // -250001
        1796: data_ff <= 24'h0271D8; // 160216
        1797: data_ff <= 24'hFE6C90; // -103280
        1798: data_ff <= 24'h00FFCC; // 65484
        1799: data_ff <= 24'hFF62D3; // -40237
        1800: data_ff <= 24'h005C76; // 23670
        1801: data_ff <= 24'hFFCC8C; // -13172
        1802: data_ff <= 24'h001AB7; // 6839
        1803: data_ff <= 24'hFFF349; // -3255
        1804: data_ff <= 24'h000568; // 1384
        1805: data_ff <= 24'hFFFE09; // -503
        1806: data_ff <= 24'h00008E; // 142
        1807: data_ff <= 24'hFFFFEB; // -21
        1808: data_ff <= 24'h374735; // 3622709
        1809: data_ff <= 24'hF40D45; // -783035
        1810: data_ff <= 24'h062D1C; // 404764
        1811: data_ff <= 24'hFC3BC9; // -246839
        1812: data_ff <= 24'h0269B4; // 158132
        1813: data_ff <= 24'hFE71E3; // -101917
        1814: data_ff <= 24'h00FC67; // 64615
        1815: data_ff <= 24'hFF64E9; // -39703
        1816: data_ff <= 24'h005B3D; // 23357
        1817: data_ff <= 24'hFFCD39; // -12999
        1818: data_ff <= 24'h001A5F; // 6751
        1819: data_ff <= 24'hFFF372; // -3214
        1820: data_ff <= 24'h000557; // 1367
        1821: data_ff <= 24'hFFFE0E; // -498
        1822: data_ff <= 24'h00008D; // 141
        1823: data_ff <= 24'hFFFFEB; // -21
        1824: data_ff <= 24'h37A0CA; // 3645642
        1825: data_ff <= 24'hF42D4A; // -774838
        1826: data_ff <= 24'h061953; // 399699
        1827: data_ff <= 24'hFC4896; // -243562
        1828: data_ff <= 24'h026145; // 155973
        1829: data_ff <= 24'hFE7766; // -100506
        1830: data_ff <= 24'h00F8E3; // 63715
        1831: data_ff <= 24'hFF6713; // -39149
        1832: data_ff <= 24'h0059F9; // 23033
        1833: data_ff <= 24'hFFCDEB; // -12821
        1834: data_ff <= 24'h001A04; // 6660
        1835: data_ff <= 24'hFFF39C; // -3172
        1836: data_ff <= 24'h000546; // 1350
        1837: data_ff <= 24'hFFFE14; // -492
        1838: data_ff <= 24'h00008B; // 139
        1839: data_ff <= 24'hFFFFEB; // -21
        1840: data_ff <= 24'h37F8C0; // 3668160
        1841: data_ff <= 24'hF44ED4; // -766252
        1842: data_ff <= 24'h0604CC; // 394444
        1843: data_ff <= 24'hFC55D5; // -240171
        1844: data_ff <= 24'h02588F; // 153743
        1845: data_ff <= 24'hFE7D18; // -99048
        1846: data_ff <= 24'h00F541; // 62785
        1847: data_ff <= 24'hFF694F; // -38577
        1848: data_ff <= 24'h0058A9; // 22697
        1849: data_ff <= 24'hFFCEA5; // -12635
        1850: data_ff <= 24'h0019A5; // 6565
        1851: data_ff <= 24'hFFF3C9; // -3127
        1852: data_ff <= 24'h000534; // 1332
        1853: data_ff <= 24'hFFFE1A; // -486
        1854: data_ff <= 24'h00008A; // 138
        1855: data_ff <= 24'hFFFFEB; // -21
        1856: data_ff <= 24'h384F10; // 3690256
        1857: data_ff <= 24'hF471E5; // -757275
        1858: data_ff <= 24'h05EF87; // 388999
        1859: data_ff <= 24'hFC6385; // -236667
        1860: data_ff <= 24'h024F8F; // 151439
        1861: data_ff <= 24'hFE82F8; // -97544
        1862: data_ff <= 24'h00F180; // 61824
        1863: data_ff <= 24'hFF6B9F; // -37985
        1864: data_ff <= 24'h00574E; // 22350
        1865: data_ff <= 24'hFFCF64; // -12444
        1866: data_ff <= 24'h001943; // 6467
        1867: data_ff <= 24'hFFF3F6; // -3082
        1868: data_ff <= 24'h000521; // 1313
        1869: data_ff <= 24'hFFFE21; // -479
        1870: data_ff <= 24'h000088; // 136
        1871: data_ff <= 24'hFFFFEB; // -21
        1872: data_ff <= 24'h38A3B7; // 3711927
        1873: data_ff <= 24'hF4967C; // -747908
        1874: data_ff <= 24'h05D984; // 383364
        1875: data_ff <= 24'hFC71A6; // -233050
        1876: data_ff <= 24'h024648; // 149064
        1877: data_ff <= 24'hFE8908; // -95992
        1878: data_ff <= 24'h00EDA2; // 60834
        1879: data_ff <= 24'hFF6E01; // -37375
        1880: data_ff <= 24'h0055E8; // 21992
        1881: data_ff <= 24'hFFD02B; // -12245
        1882: data_ff <= 24'h0018DD; // 6365
        1883: data_ff <= 24'hFFF426; // -3034
        1884: data_ff <= 24'h00050D; // 1293
        1885: data_ff <= 24'hFFFE27; // -473
        1886: data_ff <= 24'h000086; // 134
        1887: data_ff <= 24'hFFFFEB; // -21
        1888: data_ff <= 24'h38F6AE; // 3733166
        1889: data_ff <= 24'hF4BC9C; // -738148
        1890: data_ff <= 24'h05C2C6; // 377542
        1891: data_ff <= 24'hFC8037; // -229321
        1892: data_ff <= 24'h023CBA; // 146618
        1893: data_ff <= 24'hFE8F45; // -94395
        1894: data_ff <= 24'h00E9A5; // 59813
        1895: data_ff <= 24'hFF7075; // -36747
        1896: data_ff <= 24'h005476; // 21622
        1897: data_ff <= 24'hFFD0F7; // -12041
        1898: data_ff <= 24'h001874; // 6260
        1899: data_ff <= 24'hFFF457; // -2985
        1900: data_ff <= 24'h0004F9; // 1273
        1901: data_ff <= 24'hFFFE2F; // -465
        1902: data_ff <= 24'h000085; // 133
        1903: data_ff <= 24'hFFFFEB; // -21
        1904: data_ff <= 24'h3947F1; // 3753969
        1905: data_ff <= 24'hF4E446; // -727994
        1906: data_ff <= 24'h05AB4C; // 371532
        1907: data_ff <= 24'hFC8F36; // -225482
        1908: data_ff <= 24'h0232E5; // 144101
        1909: data_ff <= 24'hFE95B1; // -92751
        1910: data_ff <= 24'h00E58C; // 58764
        1911: data_ff <= 24'hFF72FD; // -36099
        1912: data_ff <= 24'h0052FA; // 21242
        1913: data_ff <= 24'hFFD1CA; // -11830
        1914: data_ff <= 24'h001807; // 6151
        1915: data_ff <= 24'hFFF48A; // -2934
        1916: data_ff <= 24'h0004E4; // 1252
        1917: data_ff <= 24'hFFFE36; // -458
        1918: data_ff <= 24'h000083; // 131
        1919: data_ff <= 24'hFFFFEC; // -20
        1920: data_ff <= 24'h39977C; // 3774332
        1921: data_ff <= 24'hF50D79; // -717447
        1922: data_ff <= 24'h059318; // 365336
        1923: data_ff <= 24'hFC9EA4; // -221532
        1924: data_ff <= 24'h0228CA; // 141514
        1925: data_ff <= 24'hFE9C4A; // -91062
        1926: data_ff <= 24'h00E155; // 57685
        1927: data_ff <= 24'hFF7596; // -35434
        1928: data_ff <= 24'h005172; // 20850
        1929: data_ff <= 24'hFFD2A4; // -11612
        1930: data_ff <= 24'h001797; // 6039
        1931: data_ff <= 24'hFFF4BF; // -2881
        1932: data_ff <= 24'h0004CE; // 1230
        1933: data_ff <= 24'hFFFE3E; // -450
        1934: data_ff <= 24'h000081; // 129
        1935: data_ff <= 24'hFFFFEC; // -20
        1936: data_ff <= 24'h39E548; // 3794248
        1937: data_ff <= 24'hF53836; // -706506
        1938: data_ff <= 24'h057A2A; // 358954
        1939: data_ff <= 24'hFCAE7F; // -217473
        1940: data_ff <= 24'h021E69; // 138857
        1941: data_ff <= 24'hFEA310; // -89328
        1942: data_ff <= 24'h00DD01; // 56577
        1943: data_ff <= 24'hFF7842; // -34750
        1944: data_ff <= 24'h004FDF; // 20447
        1945: data_ff <= 24'hFFD384; // -11388
        1946: data_ff <= 24'h001723; // 5923
        1947: data_ff <= 24'hFFF4F5; // -2827
        1948: data_ff <= 24'h0004B7; // 1207
        1949: data_ff <= 24'hFFFE45; // -443
        1950: data_ff <= 24'h00007F; // 127
        1951: data_ff <= 24'hFFFFEC; // -20
        1952: data_ff <= 24'h3A3152; // 3813714
        1953: data_ff <= 24'hF5647E; // -695170
        1954: data_ff <= 24'h056085; // 352389
        1955: data_ff <= 24'hFCBEC6; // -213306
        1956: data_ff <= 24'h0213C4; // 136132
        1957: data_ff <= 24'hFEAA03; // -87549
        1958: data_ff <= 24'h00D890; // 55440
        1959: data_ff <= 24'hFF7B00; // -34048
        1960: data_ff <= 24'h004E41; // 20033
        1961: data_ff <= 24'hFFD46A; // -11158
        1962: data_ff <= 24'h0016AC; // 5804
        1963: data_ff <= 24'hFFF52D; // -2771
        1964: data_ff <= 24'h0004A0; // 1184
        1965: data_ff <= 24'hFFFE4E; // -434
        1966: data_ff <= 24'h00007D; // 125
        1967: data_ff <= 24'hFFFFEC; // -20
        1968: data_ff <= 24'h3A7B95; // 3832725
        1969: data_ff <= 24'hF59252; // -683438
        1970: data_ff <= 24'h054628; // 345640
        1971: data_ff <= 24'hFCCF78; // -209032
        1972: data_ff <= 24'h0208DB; // 133339
        1973: data_ff <= 24'hFEB121; // -85727
        1974: data_ff <= 24'h00D403; // 54275
        1975: data_ff <= 24'hFF7DD0; // -33328
        1976: data_ff <= 24'h004C99; // 19609
        1977: data_ff <= 24'hFFD556; // -10922
        1978: data_ff <= 24'h001632; // 5682
        1979: data_ff <= 24'hFFF567; // -2713
        1980: data_ff <= 24'h000488; // 1160
        1981: data_ff <= 24'hFFFE56; // -426
        1982: data_ff <= 24'h00007A; // 122
        1983: data_ff <= 24'hFFFFEC; // -20
        1984: data_ff <= 24'h3AC40D; // 3851277
        1985: data_ff <= 24'hF5C1B1; // -671311
        1986: data_ff <= 24'h052B16; // 338710
        1987: data_ff <= 24'hFCE095; // -204651
        1988: data_ff <= 24'h01FDAE; // 130478
        1989: data_ff <= 24'hFEB86C; // -83860
        1990: data_ff <= 24'h00CF5A; // 53082
        1991: data_ff <= 24'hFF80B1; // -32591
        1992: data_ff <= 24'h004AE5; // 19173
        1993: data_ff <= 24'hFFD649; // -10679
        1994: data_ff <= 24'h0015B4; // 5556
        1995: data_ff <= 24'hFFF5A3; // -2653
        1996: data_ff <= 24'h00046F; // 1135
        1997: data_ff <= 24'hFFFE5F; // -417
        1998: data_ff <= 24'h000078; // 120
        1999: data_ff <= 24'hFFFFED; // -19
        2000: data_ff <= 24'h3B0AB4; // 3869364
        2001: data_ff <= 24'hF5F29C; // -658788
        2002: data_ff <= 24'h050F50; // 331600
        2003: data_ff <= 24'hFCF21B; // -200165
        2004: data_ff <= 24'h01F23E; // 127550
        2005: data_ff <= 24'hFEBFE2; // -81950
        2006: data_ff <= 24'h00CA94; // 51860
        2007: data_ff <= 24'hFF83A4; // -31836
        2008: data_ff <= 24'h004927; // 18727
        2009: data_ff <= 24'hFFD741; // -10431
        2010: data_ff <= 24'h001533; // 5427
        2011: data_ff <= 24'hFFF5E0; // -2592
        2012: data_ff <= 24'h000455; // 1109
        2013: data_ff <= 24'hFFFE68; // -408
        2014: data_ff <= 24'h000075; // 117
        2015: data_ff <= 24'hFFFFED; // -19
        2016: data_ff <= 24'h3B4F88; // 3886984
        2017: data_ff <= 24'hF62513; // -645869
        2018: data_ff <= 24'h04F2D7; // 324311
        2019: data_ff <= 24'hFD0409; // -195575
        2020: data_ff <= 24'h01E68D; // 124557
        2021: data_ff <= 24'hFEC782; // -79998
        2022: data_ff <= 24'h00C5B4; // 50612
        2023: data_ff <= 24'hFF86A8; // -31064
        2024: data_ff <= 24'h00475F; // 18271
        2025: data_ff <= 24'hFFD840; // -10176
        2026: data_ff <= 24'h0014AF; // 5295
        2027: data_ff <= 24'hFFF61F; // -2529
        2028: data_ff <= 24'h00043A; // 1082
        2029: data_ff <= 24'hFFFE72; // -398
        2030: data_ff <= 24'h000073; // 115
        2031: data_ff <= 24'hFFFFED; // -19
        2032: data_ff <= 24'h3B9283; // 3904131
        2033: data_ff <= 24'hF65915; // -632555
        2034: data_ff <= 24'h04D5AD; // 316845
        2035: data_ff <= 24'hFD165D; // -190883
        2036: data_ff <= 24'h01DA9B; // 121499
        2037: data_ff <= 24'hFECF4C; // -78004
        2038: data_ff <= 24'h00C0B8; // 49336
        2039: data_ff <= 24'hFF89BE; // -30274
        2040: data_ff <= 24'h00458C; // 17804
        2041: data_ff <= 24'hFFD945; // -9915
        2042: data_ff <= 24'h001427; // 5159
        2043: data_ff <= 24'hFFF65F; // -2465
        2044: data_ff <= 24'h00041F; // 1055
        2045: data_ff <= 24'hFFFE7C; // -388
        2046: data_ff <= 24'h000070; // 112
        2047: data_ff <= 24'hFFFFEE; // -18
        2048: data_ff <= 24'h3BD3A2; // 3920802
        2049: data_ff <= 24'hF68EA4; // -618844
        2050: data_ff <= 24'h04B7D3; // 309203
        2051: data_ff <= 24'hFD2918; // -186088
        2052: data_ff <= 24'h01CE68; // 118376
        2053: data_ff <= 24'hFED740; // -75968
        2054: data_ff <= 24'h00BBA1; // 48033
        2055: data_ff <= 24'hFF8CE4; // -29468
        2056: data_ff <= 24'h0043AF; // 17327
        2057: data_ff <= 24'hFFDA50; // -9648
        2058: data_ff <= 24'h00139C; // 5020
        2059: data_ff <= 24'hFFF6A1; // -2399
        2060: data_ff <= 24'h000403; // 1027
        2061: data_ff <= 24'hFFFE86; // -378
        2062: data_ff <= 24'h00006D; // 109
        2063: data_ff <= 24'hFFFFEE; // -18
        2064: data_ff <= 24'h3C12E1; // 3936993
        2065: data_ff <= 24'hF6C5BD; // -604739
        2066: data_ff <= 24'h04994B; // 301387
        2067: data_ff <= 24'hFD3C36; // -181194
        2068: data_ff <= 24'h01C1F6; // 115190
        2069: data_ff <= 24'hFEDF5E; // -73890
        2070: data_ff <= 24'h00B670; // 46704
        2071: data_ff <= 24'hFF901B; // -28645
        2072: data_ff <= 24'h0041C7; // 16839
        2073: data_ff <= 24'hFFDB60; // -9376
        2074: data_ff <= 24'h00130E; // 4878
        2075: data_ff <= 24'hFFF6E5; // -2331
        2076: data_ff <= 24'h0003E6; // 998
        2077: data_ff <= 24'hFFFE90; // -368
        2078: data_ff <= 24'h00006B; // 107
        2079: data_ff <= 24'hFFFFEE; // -18
        2080: data_ff <= 24'h3C503C; // 3952700
        2081: data_ff <= 24'hF6FE62; // -590238
        2082: data_ff <= 24'h047A17; // 293399
        2083: data_ff <= 24'hFD4FB8; // -176200
        2084: data_ff <= 24'h01B546; // 111942
        2085: data_ff <= 24'hFEE7A3; // -71773
        2086: data_ff <= 24'h00B125; // 45349
        2087: data_ff <= 24'hFF9362; // -27806
        2088: data_ff <= 24'h003FD6; // 16342
        2089: data_ff <= 24'hFFDC77; // -9097
        2090: data_ff <= 24'h00127C; // 4732
        2091: data_ff <= 24'hFFF72B; // -2261
        2092: data_ff <= 24'h0003C8; // 968
        2093: data_ff <= 24'hFFFE9B; // -357
        2094: data_ff <= 24'h000068; // 104
        2095: data_ff <= 24'hFFFFEF; // -17
        2096: data_ff <= 24'h3C8BAF; // 3967919
        2097: data_ff <= 24'hF73891; // -575343
        2098: data_ff <= 24'h045A39; // 285241
        2099: data_ff <= 24'hFD639B; // -171109
        2100: data_ff <= 24'h01A859; // 108633
        2101: data_ff <= 24'hFEF010; // -69616
        2102: data_ff <= 24'h00ABC0; // 43968
        2103: data_ff <= 24'hFF96BA; // -26950
        2104: data_ff <= 24'h003DDB; // 15835
        2105: data_ff <= 24'hFFDD93; // -8813
        2106: data_ff <= 24'h0011E8; // 4584
        2107: data_ff <= 24'hFFF772; // -2190
        2108: data_ff <= 24'h0003AA; // 938
        2109: data_ff <= 24'hFFFEA6; // -346
        2110: data_ff <= 24'h000065; // 101
        2111: data_ff <= 24'hFFFFEF; // -17
        2112: data_ff <= 24'h3CC537; // 3982647
        2113: data_ff <= 24'hF7744A; // -560054
        2114: data_ff <= 24'h0439B2; // 276914
        2115: data_ff <= 24'hFD77DF; // -165921
        2116: data_ff <= 24'h019B2E; // 105262
        2117: data_ff <= 24'hFEF8A5; // -67419
        2118: data_ff <= 24'h00A642; // 42562
        2119: data_ff <= 24'hFF9A22; // -26078
        2120: data_ff <= 24'h003BD6; // 15318
        2121: data_ff <= 24'hFFDEB5; // -8523
        2122: data_ff <= 24'h001150; // 4432
        2123: data_ff <= 24'hFFF7BA; // -2118
        2124: data_ff <= 24'h00038B; // 907
        2125: data_ff <= 24'hFFFEB1; // -335
        2126: data_ff <= 24'h000061; // 97
        2127: data_ff <= 24'hFFFFF0; // -16
        2128: data_ff <= 24'h3CFCD0; // 3996880
        2129: data_ff <= 24'hF7B18D; // -544371
        2130: data_ff <= 24'h041885; // 268421
        2131: data_ff <= 24'hFD8C81; // -160639
        2132: data_ff <= 24'h018DC9; // 101833
        2133: data_ff <= 24'hFF0160; // -65184
        2134: data_ff <= 24'h00A0AB; // 41131
        2135: data_ff <= 24'hFF9D99; // -25191
        2136: data_ff <= 24'h0039C7; // 14791
        2137: data_ff <= 24'hFFDFDD; // -8227
        2138: data_ff <= 24'h0010B5; // 4277
        2139: data_ff <= 24'hFFF805; // -2043
        2140: data_ff <= 24'h00036B; // 875
        2141: data_ff <= 24'hFFFEBD; // -323
        2142: data_ff <= 24'h00005E; // 94
        2143: data_ff <= 24'hFFFFF0; // -16
        2144: data_ff <= 24'h3D3277; // 4010615
        2145: data_ff <= 24'hF7F058; // -528296
        2146: data_ff <= 24'h03F6B3; // 259763
        2147: data_ff <= 24'hFDA181; // -155263
        2148: data_ff <= 24'h018029; // 98345
        2149: data_ff <= 24'hFF0A41; // -62911
        2150: data_ff <= 24'h009AFB; // 39675
        2151: data_ff <= 24'hFFA120; // -24288
        2152: data_ff <= 24'h0037AF; // 14255
        2153: data_ff <= 24'hFFE10A; // -7926
        2154: data_ff <= 24'h001018; // 4120
        2155: data_ff <= 24'hFFF850; // -1968
        2156: data_ff <= 24'h00034B; // 843
        2157: data_ff <= 24'hFFFEC9; // -311
        2158: data_ff <= 24'h00005B; // 91
        2159: data_ff <= 24'hFFFFF1; // -15
        2160: data_ff <= 24'h3D6629; // 4023849
        2161: data_ff <= 24'hF830AA; // -511830
        2162: data_ff <= 24'h03D43E; // 250942
        2163: data_ff <= 24'hFDB6DC; // -149796
        2164: data_ff <= 24'h01724F; // 94799
        2165: data_ff <= 24'hFF1346; // -60602
        2166: data_ff <= 24'h009534; // 38196
        2167: data_ff <= 24'hFFA4B7; // -23369
        2168: data_ff <= 24'h00358D; // 13709
        2169: data_ff <= 24'hFFE23D; // -7619
        2170: data_ff <= 24'h000F77; // 3959
        2171: data_ff <= 24'hFFF89E; // -1890
        2172: data_ff <= 24'h00032A; // 810
        2173: data_ff <= 24'hFFFED5; // -299
        2174: data_ff <= 24'h000057; // 87
        2175: data_ff <= 24'hFFFFF1; // -15
        2176: data_ff <= 24'h3D97E2; // 4036578
        2177: data_ff <= 24'hF87283; // -494973
        2178: data_ff <= 24'h03B12A; // 241962
        2179: data_ff <= 24'hFDCC92; // -144238
        2180: data_ff <= 24'h01643D; // 91197
        2181: data_ff <= 24'hFF1C71; // -58255
        2182: data_ff <= 24'h008F55; // 36693
        2183: data_ff <= 24'hFFA85C; // -22436
        2184: data_ff <= 24'h003362; // 13154
        2185: data_ff <= 24'hFFE375; // -7307
        2186: data_ff <= 24'h000ED3; // 3795
        2187: data_ff <= 24'hFFF8ED; // -1811
        2188: data_ff <= 24'h000308; // 776
        2189: data_ff <= 24'hFFFEE2; // -286
        2190: data_ff <= 24'h000054; // 84
        2191: data_ff <= 24'hFFFFF2; // -14
        2192: data_ff <= 24'h3DC7A0; // 4048800
        2193: data_ff <= 24'hF8B5E1; // -477727
        2194: data_ff <= 24'h038D77; // 232823
        2195: data_ff <= 24'hFDE2A0; // -138592
        2196: data_ff <= 24'h0155F4; // 87540
        2197: data_ff <= 24'hFF25BF; // -55873
        2198: data_ff <= 24'h00895F; // 35167
        2199: data_ff <= 24'hFFAC10; // -21488
        2200: data_ff <= 24'h00312F; // 12591
        2201: data_ff <= 24'hFFE4B2; // -6990
        2202: data_ff <= 24'h000E2C; // 3628
        2203: data_ff <= 24'hFFF93D; // -1731
        2204: data_ff <= 24'h0002E5; // 741
        2205: data_ff <= 24'hFFFEEE; // -274
        2206: data_ff <= 24'h000050; // 80
        2207: data_ff <= 24'hFFFFF2; // -14
        2208: data_ff <= 24'h3DF55F; // 4060511
        2209: data_ff <= 24'hF8FAC4; // -460092
        2210: data_ff <= 24'h036929; // 223529
        2211: data_ff <= 24'hFDF905; // -132859
        2212: data_ff <= 24'h014775; // 83829
        2213: data_ff <= 24'hFF2F30; // -53456
        2214: data_ff <= 24'h008352; // 33618
        2215: data_ff <= 24'hFFAFD2; // -20526
        2216: data_ff <= 24'h002EF2; // 12018
        2217: data_ff <= 24'hFFE5F4; // -6668
        2218: data_ff <= 24'h000D83; // 3459
        2219: data_ff <= 24'hFFF98F; // -1649
        2220: data_ff <= 24'h0002C2; // 706
        2221: data_ff <= 24'hFFFEFC; // -260
        2222: data_ff <= 24'h00004C; // 76
        2223: data_ff <= 24'hFFFFF3; // -13
        2224: data_ff <= 24'h3E211D; // 4071709
        2225: data_ff <= 24'hF9412A; // -442070
        2226: data_ff <= 24'h034442; // 214082
        2227: data_ff <= 24'hFE0FBF; // -127041
        2228: data_ff <= 24'h0138C0; // 80064
        2229: data_ff <= 24'hFF38C3; // -51005
        2230: data_ff <= 24'h007D2F; // 32047
        2231: data_ff <= 24'hFFB3A2; // -19550
        2232: data_ff <= 24'h002CAD; // 11437
        2233: data_ff <= 24'hFFE73C; // -6340
        2234: data_ff <= 24'h000CD6; // 3286
        2235: data_ff <= 24'hFFF9E2; // -1566
        2236: data_ff <= 24'h00029E; // 670
        2237: data_ff <= 24'hFFFF09; // -247
        2238: data_ff <= 24'h000048; // 72
        2239: data_ff <= 24'hFFFFF4; // -12
        2240: data_ff <= 24'h3E4AD7; // 4082391
        2241: data_ff <= 24'hF98910; // -423664
        2242: data_ff <= 24'h031EC4; // 204484
        2243: data_ff <= 24'hFE26CC; // -121140
        2244: data_ff <= 24'h0129D8; // 76248
        2245: data_ff <= 24'hFF4278; // -48520
        2246: data_ff <= 24'h0076F6; // 30454
        2247: data_ff <= 24'hFFB780; // -18560
        2248: data_ff <= 24'h002A5F; // 10847
        2249: data_ff <= 24'hFFE889; // -6007
        2250: data_ff <= 24'h000C27; // 3111
        2251: data_ff <= 24'hFFFA37; // -1481
        2252: data_ff <= 24'h000279; // 633
        2253: data_ff <= 24'hFFFF17; // -233
        2254: data_ff <= 24'h000044; // 68
        2255: data_ff <= 24'hFFFFF4; // -12
        2256: data_ff <= 24'h3E728B; // 4092555
        2257: data_ff <= 24'hF9D277; // -404873
        2258: data_ff <= 24'h02F8B1; // 194737
        2259: data_ff <= 24'hFE3E2B; // -115157
        2260: data_ff <= 24'h011ABD; // 72381
        2261: data_ff <= 24'hFF4C4E; // -46002
        2262: data_ff <= 24'h0070A8; // 28840
        2263: data_ff <= 24'hFFBB6C; // -17556
        2264: data_ff <= 24'h002809; // 10249
        2265: data_ff <= 24'hFFE9DA; // -5670
        2266: data_ff <= 24'h000B75; // 2933
        2267: data_ff <= 24'hFFFA8D; // -1395
        2268: data_ff <= 24'h000253; // 595
        2269: data_ff <= 24'hFFFF25; // -219
        2270: data_ff <= 24'h000040; // 64
        2271: data_ff <= 24'hFFFFF5; // -11
        2272: data_ff <= 24'h3E9836; // 4102198
        2273: data_ff <= 24'hFA1D5B; // -385701
        2274: data_ff <= 24'h02D20E; // 184846
        2275: data_ff <= 24'hFE55DA; // -109094
        2276: data_ff <= 24'h010B71; // 68465
        2277: data_ff <= 24'hFF5643; // -43453
        2278: data_ff <= 24'h006A46; // 27206
        2279: data_ff <= 24'hFFBF65; // -16539
        2280: data_ff <= 24'h0025AB; // 9643
        2281: data_ff <= 24'hFFEB31; // -5327
        2282: data_ff <= 24'h000AC0; // 2752
        2283: data_ff <= 24'hFFFAE5; // -1307
        2284: data_ff <= 24'h00022D; // 557
        2285: data_ff <= 24'hFFFF33; // -205
        2286: data_ff <= 24'h00003C; // 60
        2287: data_ff <= 24'hFFFFF6; // -10
        2288: data_ff <= 24'h3EBBD6; // 4111318
        2289: data_ff <= 24'hFA69BC; // -366148
        2290: data_ff <= 24'h02AADB; // 174811
        2291: data_ff <= 24'hFE6DD7; // -102953
        2292: data_ff <= 24'h00FBF5; // 64501
        2293: data_ff <= 24'hFF6057; // -40873
        2294: data_ff <= 24'h0063CF; // 25551
        2295: data_ff <= 24'hFFC36A; // -15510
        2296: data_ff <= 24'h002344; // 9028
        2297: data_ff <= 24'hFFEC8C; // -4980
        2298: data_ff <= 24'h000A09; // 2569
        2299: data_ff <= 24'hFFFB3E; // -1218
        2300: data_ff <= 24'h000207; // 519
        2301: data_ff <= 24'hFFFF41; // -191
        2302: data_ff <= 24'h000038; // 56
        2303: data_ff <= 24'hFFFFF6; // -10
        2304: data_ff <= 24'h3EDD68; // 4119912
        2305: data_ff <= 24'hFAB798; // -346216
        2306: data_ff <= 24'h02831C; // 164636
        2307: data_ff <= 24'hFE8620; // -96736
        2308: data_ff <= 24'h00EC4A; // 60490
        2309: data_ff <= 24'hFF6A89; // -38263
        2310: data_ff <= 24'h005D45; // 23877
        2311: data_ff <= 24'hFFC77C; // -14468
        2312: data_ff <= 24'h0020D6; // 8406
        2313: data_ff <= 24'hFFEDEC; // -4628
        2314: data_ff <= 24'h00094F; // 2383
        2315: data_ff <= 24'hFFFB98; // -1128
        2316: data_ff <= 24'h0001DF; // 479
        2317: data_ff <= 24'hFFFF50; // -176
        2318: data_ff <= 24'h000033; // 51
        2319: data_ff <= 24'hFFFFF7; // -9
        2320: data_ff <= 24'h3EFCEC; // 4127980
        2321: data_ff <= 24'hFB06EB; // -325909
        2322: data_ff <= 24'h025AD4; // 154324
        2323: data_ff <= 24'hFE9EB2; // -90446
        2324: data_ff <= 24'h00DC72; // 56434
        2325: data_ff <= 24'hFF74D9; // -35623
        2326: data_ff <= 24'h0056A8; // 22184
        2327: data_ff <= 24'hFFCB9A; // -13414
        2328: data_ff <= 24'h001E61; // 7777
        2329: data_ff <= 24'hFFEF50; // -4272
        2330: data_ff <= 24'h000892; // 2194
        2331: data_ff <= 24'hFFFBF4; // -1036
        2332: data_ff <= 24'h0001B7; // 439
        2333: data_ff <= 24'hFFFF5F; // -161
        2334: data_ff <= 24'h00002F; // 47
        2335: data_ff <= 24'hFFFFF8; // -8
        2336: data_ff <= 24'h3F1A5E; // 4135518
        2337: data_ff <= 24'hFB57B5; // -305227
        2338: data_ff <= 24'h023206; // 143878
        2339: data_ff <= 24'hFEB78D; // -84083
        2340: data_ff <= 24'h00CC6E; // 52334
        2341: data_ff <= 24'hFF7F45; // -32955
        2342: data_ff <= 24'h004FF8; // 20472
        2343: data_ff <= 24'hFFCFC5; // -12347
        2344: data_ff <= 24'h001BE4; // 7140
        2345: data_ff <= 24'hFFF0B8; // -3912
        2346: data_ff <= 24'h0007D3; // 2003
        2347: data_ff <= 24'hFFFC51; // -943
        2348: data_ff <= 24'h00018E; // 398
        2349: data_ff <= 24'hFFFF6F; // -145
        2350: data_ff <= 24'h00002A; // 42
        2351: data_ff <= 24'hFFFFF9; // -7
        2352: data_ff <= 24'h3F35BD; // 4142525
        2353: data_ff <= 24'hFBA9F3; // -284173
        2354: data_ff <= 24'h0208B4; // 133300
        2355: data_ff <= 24'hFED0AD; // -77651
        2356: data_ff <= 24'h00BC3E; // 48190
        2357: data_ff <= 24'hFF89CD; // -30259
        2358: data_ff <= 24'h004937; // 18743
        2359: data_ff <= 24'hFFD3FA; // -11270
        2360: data_ff <= 24'h001960; // 6496
        2361: data_ff <= 24'hFFF225; // -3547
        2362: data_ff <= 24'h000712; // 1810
        2363: data_ff <= 24'hFFFCAF; // -849
        2364: data_ff <= 24'h000165; // 357
        2365: data_ff <= 24'hFFFF7E; // -130
        2366: data_ff <= 24'h000025; // 37
        2367: data_ff <= 24'hFFFFFA; // -6
        2368: data_ff <= 24'h3F4F08; // 4149000
        2369: data_ff <= 24'hFBFDA2; // -262750
        2370: data_ff <= 24'h01DEE2; // 122594
        2371: data_ff <= 24'hFEEA12; // -71150
        2372: data_ff <= 24'h00ABE6; // 44006
        2373: data_ff <= 24'hFF946F; // -27537
        2374: data_ff <= 24'h004264; // 16996
        2375: data_ff <= 24'hFFD83B; // -10181
        2376: data_ff <= 24'h0016D5; // 5845
        2377: data_ff <= 24'hFFF396; // -3178
        2378: data_ff <= 24'h00064E; // 1614
        2379: data_ff <= 24'hFFFD0F; // -753
        2380: data_ff <= 24'h00013B; // 315
        2381: data_ff <= 24'hFFFF8E; // -114
        2382: data_ff <= 24'h000021; // 33
        2383: data_ff <= 24'hFFFFFB; // -5
        2384: data_ff <= 24'h3F663D; // 4154941
        2385: data_ff <= 24'hFC52C1; // -240959
        2386: data_ff <= 24'h01B493; // 111763
        2387: data_ff <= 24'hFF03B8; // -64584
        2388: data_ff <= 24'h009B65; // 39781
        2389: data_ff <= 24'hFF9F2B; // -24789
        2390: data_ff <= 24'h003B81; // 15233
        2391: data_ff <= 24'hFFDC86; // -9082
        2392: data_ff <= 24'h001443; // 5187
        2393: data_ff <= 24'hFFF50B; // -2805
        2394: data_ff <= 24'h000588; // 1416
        2395: data_ff <= 24'hFFFD70; // -656
        2396: data_ff <= 24'h000111; // 273
        2397: data_ff <= 24'hFFFF9E; // -98
        2398: data_ff <= 24'h00001C; // 28
        2399: data_ff <= 24'hFFFFFC; // -4
        2400: data_ff <= 24'h3F7B5A; // 4160346
        2401: data_ff <= 24'hFCA94C; // -218804
        2402: data_ff <= 24'h0189C9; // 100809
        2403: data_ff <= 24'hFF1D9D; // -57955
        2404: data_ff <= 24'h008ABE; // 35518
        2405: data_ff <= 24'hFFA9FF; // -22017
        2406: data_ff <= 24'h00348D; // 13453
        2407: data_ff <= 24'hFFE0DC; // -7972
        2408: data_ff <= 24'h0011AB; // 4523
        2409: data_ff <= 24'hFFF684; // -2428
        2410: data_ff <= 24'h0004C0; // 1216
        2411: data_ff <= 24'hFFFDD2; // -558
        2412: data_ff <= 24'h0000E6; // 230
        2413: data_ff <= 24'hFFFFAF; // -81
        2414: data_ff <= 24'h000017; // 23
        2415: data_ff <= 24'hFFFFFC; // -4
        2416: data_ff <= 24'h3F8E5E; // 4165214
        2417: data_ff <= 24'hFD0141; // -196287
        2418: data_ff <= 24'h015E89; // 89737
        2419: data_ff <= 24'hFF37C0; // -51264
        2420: data_ff <= 24'h0079F2; // 31218
        2421: data_ff <= 24'hFFB4EB; // -19221
        2422: data_ff <= 24'h002D8A; // 11658
        2423: data_ff <= 24'hFFE53C; // -6852
        2424: data_ff <= 24'h000F0D; // 3853
        2425: data_ff <= 24'hFFF801; // -2047
        2426: data_ff <= 24'h0003F5; // 1013
        2427: data_ff <= 24'hFFFE35; // -459
        2428: data_ff <= 24'h0000BA; // 186
        2429: data_ff <= 24'hFFFFBF; // -65
        2430: data_ff <= 24'h000012; // 18
        2431: data_ff <= 24'hFFFFFD; // -3
        2432: data_ff <= 24'h3F9F48; // 4169544
        2433: data_ff <= 24'hFD5A9E; // -173410
        2434: data_ff <= 24'h0132D5; // 78549
        2435: data_ff <= 24'hFF521F; // -44513
        2436: data_ff <= 24'h006902; // 26882
        2437: data_ff <= 24'hFFBFEF; // -16401
        2438: data_ff <= 24'h002678; // 9848
        2439: data_ff <= 24'hFFE9A5; // -5723
        2440: data_ff <= 24'h000C68; // 3176
        2441: data_ff <= 24'hFFF982; // -1662
        2442: data_ff <= 24'h000329; // 809
        2443: data_ff <= 24'hFFFE99; // -359
        2444: data_ff <= 24'h00008E; // 142
        2445: data_ff <= 24'hFFFFD0; // -48
        2446: data_ff <= 24'h00000C; // 12
        2447: data_ff <= 24'hFFFFFE; // -2
        2448: data_ff <= 24'h3FAE18; // 4173336
        2449: data_ff <= 24'hFDB55E; // -150178
        2450: data_ff <= 24'h0106B1; // 67249
        2451: data_ff <= 24'hFF6CB6; // -37706
        2452: data_ff <= 24'h0057F0; // 22512
        2453: data_ff <= 24'hFFCB08; // -13560
        2454: data_ff <= 24'h001F58; // 8024
        2455: data_ff <= 24'hFFEE18; // -4584
        2456: data_ff <= 24'h0009BE; // 2494
        2457: data_ff <= 24'hFFFB06; // -1274
        2458: data_ff <= 24'h00025A; // 602
        2459: data_ff <= 24'hFFFEFE; // -258
        2460: data_ff <= 24'h000061; // 97
        2461: data_ff <= 24'hFFFFE1; // -31
        2462: data_ff <= 24'h000007; // 7
        2463: data_ff <= 24'hFFFFFF; // -1
        2464: data_ff <= 24'h3FBACB; // 4176587
        2465: data_ff <= 24'hFE1180; // -126592
        2466: data_ff <= 24'h00DA20; // 55840
        2467: data_ff <= 24'hFF8783; // -30845
        2468: data_ff <= 24'h0046BE; // 18110
        2469: data_ff <= 24'hFFD635; // -10699
        2470: data_ff <= 24'h00182A; // 6186
        2471: data_ff <= 24'hFFF293; // -3437
        2472: data_ff <= 24'h00070E; // 1806
        2473: data_ff <= 24'hFFFC8D; // -883
        2474: data_ff <= 24'h000189; // 393
        2475: data_ff <= 24'hFFFF65; // -155
        2476: data_ff <= 24'h000034; // 52
        2477: data_ff <= 24'hFFFFF3; // -13
        2478: data_ff <= 24'h000002; // 2
        2479: data_ff <= 24'h000000; // 0
        2480: data_ff <= 24'h3FC561; // 4179297
        2481: data_ff <= 24'hFE6F00; // -102656
        2482: data_ff <= 24'h00AD25; // 44325
        2483: data_ff <= 24'hFFA285; // -23931
        2484: data_ff <= 24'h00356C; // 13676
        2485: data_ff <= 24'hFFE177; // -7817
        2486: data_ff <= 24'h0010F0; // 4336
        2487: data_ff <= 24'hFFF717; // -2281
        2488: data_ff <= 24'h000459; // 1113
        2489: data_ff <= 24'hFFFE18; // -488
        2490: data_ff <= 24'h0000B7; // 183
        2491: data_ff <= 24'hFFFFCC; // -52
        2492: data_ff <= 24'h000006; // 6
        2493: data_ff <= 24'h000004; // 4
        2494: data_ff <= 24'hFFFFFD; // -3
        2495: data_ff <= 24'h000001; // 1
        2496: data_ff <= 24'h3FCDDB; // 4181467
        2497: data_ff <= 24'hFECDDB; // -78373
        2498: data_ff <= 24'h007FC5; // 32709
        2499: data_ff <= 24'hFFBDB9; // -16967
        2500: data_ff <= 24'h0023FD; // 9213
        2501: data_ff <= 24'hFFECCB; // -4917
        2502: data_ff <= 24'h0009A9; // 2473
        2503: data_ff <= 24'hFFFBA3; // -1117
        2504: data_ff <= 24'h00019E; // 414
        2505: data_ff <= 24'hFFFFA6; // -90
        2506: data_ff <= 24'hFFFFE3; // -29
        2507: data_ff <= 24'h000034; // 52
        2508: data_ff <= 24'hFFFFD8; // -40
        2509: data_ff <= 24'h000015; // 21
        2510: data_ff <= 24'hFFFFF8; // -8
        2511: data_ff <= 24'h000002; // 2
        2512: data_ff <= 24'h3FD436; // 4183094
        2513: data_ff <= 24'hFF2E0E; // -53746
        2514: data_ff <= 24'h005203; // 20995
        2515: data_ff <= 24'hFFD91D; // -9955
        2516: data_ff <= 24'h001273; // 4723
        2517: data_ff <= 24'hFFF831; // -1999
        2518: data_ff <= 24'h000256; // 598
        2519: data_ff <= 24'h000035; // 53
        2520: data_ff <= 24'hFFFEE0; // -288
        2521: data_ff <= 24'h000135; // 309
        2522: data_ff <= 24'hFFFF0D; // -243
        2523: data_ff <= 24'h00009D; // 157
        2524: data_ff <= 24'hFFFFAA; // -86
        2525: data_ff <= 24'h000027; // 39
        2526: data_ff <= 24'hFFFFF2; // -14
        2527: data_ff <= 24'h000003; // 3
        2528: data_ff <= 24'h3FD873; // 4184179
        2529: data_ff <= 24'hFF8F95; // -28779
        2530: data_ff <= 24'h0023E3; // 9187
        2531: data_ff <= 24'hFFF4AD; // -2899
        2532: data_ff <= 24'h0000CD; // 205
        2533: data_ff <= 24'h0003A7; // 935
        2534: data_ff <= 24'hFFFAFA; // -1286
        2535: data_ff <= 24'h0004CF; // 1231
        2536: data_ff <= 24'hFFFC1C; // -996
        2537: data_ff <= 24'h0002C9; // 713
        2538: data_ff <= 24'hFFFE35; // -459
        2539: data_ff <= 24'h000108; // 264
        2540: data_ff <= 24'hFFFF7A; // -134
        2541: data_ff <= 24'h00003A; // 58
        2542: data_ff <= 24'hFFFFEC; // -20
        2543: data_ff <= 24'h000004; // 4
        2544: data_ff <= 24'h3FDA92; // 4184722
        2545: data_ff <= 24'hFFF26C; // -3476
        2546: data_ff <= 24'hFFF568; // -2712
        2547: data_ff <= 24'h001067; // 4199
        2548: data_ff <= 24'hFFEF11; // -4335
        2549: data_ff <= 24'h000F2D; // 3885
        2550: data_ff <= 24'hFFF392; // -3182
        2551: data_ff <= 24'h000971; // 2417
        2552: data_ff <= 24'hFFF954; // -1708
        2553: data_ff <= 24'h000460; // 1120
        2554: data_ff <= 24'hFFFD5C; // -676
        2555: data_ff <= 24'h000173; // 371
        2556: data_ff <= 24'hFFFF4A; // -182
        2557: data_ff <= 24'h00004C; // 76
        2558: data_ff <= 24'hFFFFE6; // -26
        2559: data_ff <= 24'h000005; // 5

        default: data_ff <= 0;
    endcase
end
endmodule
