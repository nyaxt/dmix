module rom_firbank_441_480(
    input clk,
    input [11:0] addr,
    output [15:0] data);
reg [15:0] data_ff;
assign data = data_ff;
always @(posedge clk) begin
    case(addr)
        0: data_ff <= 16'd6;
        1: data_ff <= -16'd13;
        2: data_ff <= 16'd20;
        3: data_ff <= -16'd26;
        4: data_ff <= 16'd29;
        5: data_ff <= -16'd20;
        6: data_ff <= -16'd26;
        7: data_ff <= 16'd32717;
        8: data_ff <= 16'd171;
        9: data_ff <= -16'd109;
        10: data_ff <= 16'd78;
        11: data_ff <= -16'd55;
        12: data_ff <= 16'd36;
        13: data_ff <= -16'd21;
        14: data_ff <= 16'd10;
        15: data_ff <= -16'd3;
        16: data_ff <= 16'd3;
        17: data_ff <= -16'd5;
        18: data_ff <= 16'd4;
        19: data_ff <= 16'd1;
        20: data_ff <= -16'd20;
        21: data_ff <= 16'd68;
        22: data_ff <= -16'd222;
        23: data_ff <= 16'd32712;
        24: data_ff <= 16'd371;
        25: data_ff <= -16'd198;
        26: data_ff <= 16'd128;
        27: data_ff <= -16'd83;
        28: data_ff <= 16'd52;
        29: data_ff <= -16'd29;
        30: data_ff <= 16'd13;
        31: data_ff <= -16'd4;
        32: data_ff <= 16'd0;
        33: data_ff <= 16'd2;
        34: data_ff <= -16'd10;
        35: data_ff <= 16'd29;
        36: data_ff <= -16'd68;
        37: data_ff <= 16'd155;
        38: data_ff <= -16'd414;
        39: data_ff <= 16'd32704;
        40: data_ff <= 16'd574;
        41: data_ff <= -16'd289;
        42: data_ff <= 16'd178;
        43: data_ff <= -16'd112;
        44: data_ff <= 16'd67;
        45: data_ff <= -16'd37;
        46: data_ff <= 16'd16;
        47: data_ff <= -16'd5;
        48: data_ff <= -16'd3;
        49: data_ff <= 16'd10;
        50: data_ff <= -16'd25;
        51: data_ff <= 16'd57;
        52: data_ff <= -16'd117;
        53: data_ff <= 16'd242;
        54: data_ff <= -16'd604;
        55: data_ff <= 16'd32691;
        56: data_ff <= 16'd780;
        57: data_ff <= -16'd380;
        58: data_ff <= 16'd228;
        59: data_ff <= -16'd141;
        60: data_ff <= 16'd83;
        61: data_ff <= -16'd45;
        62: data_ff <= 16'd20;
        63: data_ff <= -16'd6;
        64: data_ff <= -16'd6;
        65: data_ff <= 16'd17;
        66: data_ff <= -16'd41;
        67: data_ff <= 16'd84;
        68: data_ff <= -16'd165;
        69: data_ff <= 16'd328;
        70: data_ff <= -16'd791;
        71: data_ff <= 16'd32674;
        72: data_ff <= 16'd988;
        73: data_ff <= -16'd471;
        74: data_ff <= 16'd279;
        75: data_ff <= -16'd170;
        76: data_ff <= 16'd100;
        77: data_ff <= -16'd53;
        78: data_ff <= 16'd23;
        79: data_ff <= -16'd7;
        80: data_ff <= -16'd9;
        81: data_ff <= 16'd25;
        82: data_ff <= -16'd56;
        83: data_ff <= 16'd111;
        84: data_ff <= -16'd212;
        85: data_ff <= 16'd413;
        86: data_ff <= -16'd976;
        87: data_ff <= 16'd32653;
        88: data_ff <= 16'd1199;
        89: data_ff <= -16'd563;
        90: data_ff <= 16'd330;
        91: data_ff <= -16'd199;
        92: data_ff <= 16'd116;
        93: data_ff <= -16'd61;
        94: data_ff <= 16'd27;
        95: data_ff <= -16'd8;
        96: data_ff <= -16'd12;
        97: data_ff <= 16'd32;
        98: data_ff <= -16'd71;
        99: data_ff <= 16'd139;
        100: data_ff <= -16'd260;
        101: data_ff <= 16'd498;
        102: data_ff <= -16'd1158;
        103: data_ff <= 16'd32627;
        104: data_ff <= 16'd1412;
        105: data_ff <= -16'd656;
        106: data_ff <= 16'd381;
        107: data_ff <= -16'd228;
        108: data_ff <= 16'd132;
        109: data_ff <= -16'd69;
        110: data_ff <= 16'd31;
        111: data_ff <= -16'd9;
        112: data_ff <= -16'd15;
        113: data_ff <= 16'd40;
        114: data_ff <= -16'd85;
        115: data_ff <= 16'd165;
        116: data_ff <= -16'd306;
        117: data_ff <= 16'd581;
        118: data_ff <= -16'd1337;
        119: data_ff <= 16'd32597;
        120: data_ff <= 16'd1627;
        121: data_ff <= -16'd749;
        122: data_ff <= 16'd432;
        123: data_ff <= -16'd258;
        124: data_ff <= 16'd148;
        125: data_ff <= -16'd78;
        126: data_ff <= 16'd34;
        127: data_ff <= -16'd10;
        128: data_ff <= -16'd18;
        129: data_ff <= 16'd47;
        130: data_ff <= -16'd100;
        131: data_ff <= 16'd192;
        132: data_ff <= -16'd353;
        133: data_ff <= 16'd664;
        134: data_ff <= -16'd1513;
        135: data_ff <= 16'd32563;
        136: data_ff <= 16'd1845;
        137: data_ff <= -16'd842;
        138: data_ff <= 16'd483;
        139: data_ff <= -16'd287;
        140: data_ff <= 16'd165;
        141: data_ff <= -16'd86;
        142: data_ff <= 16'd38;
        143: data_ff <= -16'd11;
        144: data_ff <= -16'd21;
        145: data_ff <= 16'd54;
        146: data_ff <= -16'd114;
        147: data_ff <= 16'd218;
        148: data_ff <= -16'd399;
        149: data_ff <= 16'd745;
        150: data_ff <= -16'd1686;
        151: data_ff <= 16'd32525;
        152: data_ff <= 16'd2065;
        153: data_ff <= -16'd936;
        154: data_ff <= 16'd535;
        155: data_ff <= -16'd317;
        156: data_ff <= 16'd181;
        157: data_ff <= -16'd95;
        158: data_ff <= 16'd41;
        159: data_ff <= -16'd12;
        160: data_ff <= -16'd24;
        161: data_ff <= 16'd61;
        162: data_ff <= -16'd129;
        163: data_ff <= 16'd244;
        164: data_ff <= -16'd444;
        165: data_ff <= 16'd826;
        166: data_ff <= -16'd1856;
        167: data_ff <= 16'd32482;
        168: data_ff <= 16'd2288;
        169: data_ff <= -16'd1031;
        170: data_ff <= 16'd587;
        171: data_ff <= -16'd347;
        172: data_ff <= 16'd198;
        173: data_ff <= -16'd103;
        174: data_ff <= 16'd45;
        175: data_ff <= -16'd13;
        176: data_ff <= -16'd27;
        177: data_ff <= 16'd68;
        178: data_ff <= -16'd143;
        179: data_ff <= 16'd270;
        180: data_ff <= -16'd489;
        181: data_ff <= 16'd906;
        182: data_ff <= -16'd2024;
        183: data_ff <= 16'd32435;
        184: data_ff <= 16'd2513;
        185: data_ff <= -16'd1126;
        186: data_ff <= 16'd639;
        187: data_ff <= -16'd377;
        188: data_ff <= 16'd214;
        189: data_ff <= -16'd111;
        190: data_ff <= 16'd49;
        191: data_ff <= -16'd14;
        192: data_ff <= -16'd30;
        193: data_ff <= 16'd75;
        194: data_ff <= -16'd157;
        195: data_ff <= 16'd296;
        196: data_ff <= -16'd533;
        197: data_ff <= 16'd985;
        198: data_ff <= -16'd2189;
        199: data_ff <= 16'd32384;
        200: data_ff <= 16'd2740;
        201: data_ff <= -16'd1221;
        202: data_ff <= 16'd691;
        203: data_ff <= -16'd406;
        204: data_ff <= 16'd231;
        205: data_ff <= -16'd120;
        206: data_ff <= 16'd53;
        207: data_ff <= -16'd16;
        208: data_ff <= -16'd33;
        209: data_ff <= 16'd82;
        210: data_ff <= -16'd171;
        211: data_ff <= 16'd321;
        212: data_ff <= -16'd577;
        213: data_ff <= 16'd1062;
        214: data_ff <= -16'd2350;
        215: data_ff <= 16'd32329;
        216: data_ff <= 16'd2969;
        217: data_ff <= -16'd1316;
        218: data_ff <= 16'd743;
        219: data_ff <= -16'd436;
        220: data_ff <= 16'd248;
        221: data_ff <= -16'd129;
        222: data_ff <= 16'd56;
        223: data_ff <= -16'd17;
        224: data_ff <= -16'd35;
        225: data_ff <= 16'd89;
        226: data_ff <= -16'd184;
        227: data_ff <= 16'd346;
        228: data_ff <= -16'd620;
        229: data_ff <= 16'd1139;
        230: data_ff <= -16'd2509;
        231: data_ff <= 16'd32270;
        232: data_ff <= 16'd3201;
        233: data_ff <= -16'd1412;
        234: data_ff <= 16'd795;
        235: data_ff <= -16'd466;
        236: data_ff <= 16'd264;
        237: data_ff <= -16'd137;
        238: data_ff <= 16'd60;
        239: data_ff <= -16'd18;
        240: data_ff <= -16'd38;
        241: data_ff <= 16'd95;
        242: data_ff <= -16'd198;
        243: data_ff <= 16'd370;
        244: data_ff <= -16'd663;
        245: data_ff <= 16'd1215;
        246: data_ff <= -16'd2665;
        247: data_ff <= 16'd32206;
        248: data_ff <= 16'd3434;
        249: data_ff <= -16'd1508;
        250: data_ff <= 16'd847;
        251: data_ff <= -16'd496;
        252: data_ff <= 16'd281;
        253: data_ff <= -16'd146;
        254: data_ff <= 16'd64;
        255: data_ff <= -16'd19;
        256: data_ff <= -16'd41;
        257: data_ff <= 16'd102;
        258: data_ff <= -16'd211;
        259: data_ff <= 16'd395;
        260: data_ff <= -16'd706;
        261: data_ff <= 16'd1290;
        262: data_ff <= -16'd2818;
        263: data_ff <= 16'd32138;
        264: data_ff <= 16'd3670;
        265: data_ff <= -16'd1604;
        266: data_ff <= 16'd899;
        267: data_ff <= -16'd526;
        268: data_ff <= 16'd298;
        269: data_ff <= -16'd154;
        270: data_ff <= 16'd68;
        271: data_ff <= -16'd20;
        272: data_ff <= -16'd43;
        273: data_ff <= 16'd108;
        274: data_ff <= -16'd224;
        275: data_ff <= 16'd418;
        276: data_ff <= -16'd747;
        277: data_ff <= 16'd1363;
        278: data_ff <= -16'd2968;
        279: data_ff <= 16'd32067;
        280: data_ff <= 16'd3908;
        281: data_ff <= -16'd1700;
        282: data_ff <= 16'd952;
        283: data_ff <= -16'd556;
        284: data_ff <= 16'd314;
        285: data_ff <= -16'd163;
        286: data_ff <= 16'd72;
        287: data_ff <= -16'd22;
        288: data_ff <= -16'd46;
        289: data_ff <= 16'd115;
        290: data_ff <= -16'd237;
        291: data_ff <= 16'd442;
        292: data_ff <= -16'd788;
        293: data_ff <= 16'd1436;
        294: data_ff <= -16'd3115;
        295: data_ff <= 16'd31991;
        296: data_ff <= 16'd4147;
        297: data_ff <= -16'd1797;
        298: data_ff <= 16'd1004;
        299: data_ff <= -16'd586;
        300: data_ff <= 16'd331;
        301: data_ff <= -16'd172;
        302: data_ff <= 16'd75;
        303: data_ff <= -16'd23;
        304: data_ff <= -16'd48;
        305: data_ff <= 16'd121;
        306: data_ff <= -16'd250;
        307: data_ff <= 16'd465;
        308: data_ff <= -16'd829;
        309: data_ff <= 16'd1507;
        310: data_ff <= -16'd3259;
        311: data_ff <= 16'd31911;
        312: data_ff <= 16'd4389;
        313: data_ff <= -16'd1893;
        314: data_ff <= 16'd1056;
        315: data_ff <= -16'd616;
        316: data_ff <= 16'd348;
        317: data_ff <= -16'd180;
        318: data_ff <= 16'd79;
        319: data_ff <= -16'd24;
        320: data_ff <= -16'd51;
        321: data_ff <= 16'd127;
        322: data_ff <= -16'd262;
        323: data_ff <= 16'd488;
        324: data_ff <= -16'd869;
        325: data_ff <= 16'd1577;
        326: data_ff <= -16'd3400;
        327: data_ff <= 16'd31827;
        328: data_ff <= 16'd4633;
        329: data_ff <= -16'd1990;
        330: data_ff <= 16'd1108;
        331: data_ff <= -16'd646;
        332: data_ff <= 16'd365;
        333: data_ff <= -16'd189;
        334: data_ff <= 16'd83;
        335: data_ff <= -16'd25;
        336: data_ff <= -16'd53;
        337: data_ff <= 16'd133;
        338: data_ff <= -16'd274;
        339: data_ff <= 16'd511;
        340: data_ff <= -16'd908;
        341: data_ff <= 16'd1646;
        342: data_ff <= -16'd3538;
        343: data_ff <= 16'd31738;
        344: data_ff <= 16'd4878;
        345: data_ff <= -16'd2086;
        346: data_ff <= 16'd1161;
        347: data_ff <= -16'd676;
        348: data_ff <= 16'd381;
        349: data_ff <= -16'd198;
        350: data_ff <= 16'd87;
        351: data_ff <= -16'd27;
        352: data_ff <= -16'd55;
        353: data_ff <= 16'd139;
        354: data_ff <= -16'd286;
        355: data_ff <= 16'd533;
        356: data_ff <= -16'd947;
        357: data_ff <= 16'd1714;
        358: data_ff <= -16'd3673;
        359: data_ff <= 16'd31646;
        360: data_ff <= 16'd5125;
        361: data_ff <= -16'd2183;
        362: data_ff <= 16'd1213;
        363: data_ff <= -16'd705;
        364: data_ff <= 16'd398;
        365: data_ff <= -16'd206;
        366: data_ff <= 16'd91;
        367: data_ff <= -16'd28;
        368: data_ff <= -16'd58;
        369: data_ff <= 16'd145;
        370: data_ff <= -16'd298;
        371: data_ff <= 16'd555;
        372: data_ff <= -16'd985;
        373: data_ff <= 16'd1781;
        374: data_ff <= -16'd3805;
        375: data_ff <= 16'd31550;
        376: data_ff <= 16'd5375;
        377: data_ff <= -16'd2279;
        378: data_ff <= 16'd1264;
        379: data_ff <= -16'd735;
        380: data_ff <= 16'd415;
        381: data_ff <= -16'd215;
        382: data_ff <= 16'd95;
        383: data_ff <= -16'd29;
        384: data_ff <= -16'd60;
        385: data_ff <= 16'd150;
        386: data_ff <= -16'd310;
        387: data_ff <= 16'd576;
        388: data_ff <= -16'd1022;
        389: data_ff <= 16'd1846;
        390: data_ff <= -16'd3934;
        391: data_ff <= 16'd31450;
        392: data_ff <= 16'd5625;
        393: data_ff <= -16'd2376;
        394: data_ff <= 16'd1316;
        395: data_ff <= -16'd765;
        396: data_ff <= 16'd431;
        397: data_ff <= -16'd224;
        398: data_ff <= 16'd99;
        399: data_ff <= -16'd31;
        400: data_ff <= -16'd62;
        401: data_ff <= 16'd156;
        402: data_ff <= -16'd321;
        403: data_ff <= 16'd597;
        404: data_ff <= -16'd1059;
        405: data_ff <= 16'd1910;
        406: data_ff <= -16'd4060;
        407: data_ff <= 16'd31345;
        408: data_ff <= 16'd5878;
        409: data_ff <= -16'd2472;
        410: data_ff <= 16'd1368;
        411: data_ff <= -16'd794;
        412: data_ff <= 16'd448;
        413: data_ff <= -16'd232;
        414: data_ff <= 16'd103;
        415: data_ff <= -16'd32;
        416: data_ff <= -16'd64;
        417: data_ff <= 16'd161;
        418: data_ff <= -16'd332;
        419: data_ff <= 16'd618;
        420: data_ff <= -16'd1095;
        421: data_ff <= 16'd1973;
        422: data_ff <= -16'd4183;
        423: data_ff <= 16'd31237;
        424: data_ff <= 16'd6132;
        425: data_ff <= -16'd2568;
        426: data_ff <= 16'd1419;
        427: data_ff <= -16'd824;
        428: data_ff <= 16'd464;
        429: data_ff <= -16'd241;
        430: data_ff <= 16'd107;
        431: data_ff <= -16'd33;
        432: data_ff <= -16'd66;
        433: data_ff <= 16'd166;
        434: data_ff <= -16'd343;
        435: data_ff <= 16'd638;
        436: data_ff <= -16'd1130;
        437: data_ff <= 16'd2035;
        438: data_ff <= -16'd4302;
        439: data_ff <= 16'd31125;
        440: data_ff <= 16'd6388;
        441: data_ff <= -16'd2664;
        442: data_ff <= 16'd1471;
        443: data_ff <= -16'd853;
        444: data_ff <= 16'd481;
        445: data_ff <= -16'd249;
        446: data_ff <= 16'd110;
        447: data_ff <= -16'd35;
        448: data_ff <= -16'd68;
        449: data_ff <= 16'd172;
        450: data_ff <= -16'd354;
        451: data_ff <= 16'd658;
        452: data_ff <= -16'd1165;
        453: data_ff <= 16'd2096;
        454: data_ff <= -16'd4419;
        455: data_ff <= 16'd31009;
        456: data_ff <= 16'd6645;
        457: data_ff <= -16'd2760;
        458: data_ff <= 16'd1522;
        459: data_ff <= -16'd882;
        460: data_ff <= 16'd497;
        461: data_ff <= -16'd258;
        462: data_ff <= 16'd114;
        463: data_ff <= -16'd36;
        464: data_ff <= -16'd70;
        465: data_ff <= 16'd177;
        466: data_ff <= -16'd365;
        467: data_ff <= 16'd677;
        468: data_ff <= -16'd1199;
        469: data_ff <= 16'd2155;
        470: data_ff <= -16'd4532;
        471: data_ff <= 16'd30889;
        472: data_ff <= 16'd6904;
        473: data_ff <= -16'd2856;
        474: data_ff <= 16'd1572;
        475: data_ff <= -16'd911;
        476: data_ff <= 16'd514;
        477: data_ff <= -16'd267;
        478: data_ff <= 16'd118;
        479: data_ff <= -16'd37;
        480: data_ff <= -16'd72;
        481: data_ff <= 16'd182;
        482: data_ff <= -16'd375;
        483: data_ff <= 16'd696;
        484: data_ff <= -16'd1232;
        485: data_ff <= 16'd2213;
        486: data_ff <= -16'd4643;
        487: data_ff <= 16'd30766;
        488: data_ff <= 16'd7164;
        489: data_ff <= -16'd2951;
        490: data_ff <= 16'd1623;
        491: data_ff <= -16'd940;
        492: data_ff <= 16'd530;
        493: data_ff <= -16'd275;
        494: data_ff <= 16'd122;
        495: data_ff <= -16'd39;
        496: data_ff <= -16'd74;
        497: data_ff <= 16'd186;
        498: data_ff <= -16'd385;
        499: data_ff <= 16'd715;
        500: data_ff <= -16'd1265;
        501: data_ff <= 16'd2269;
        502: data_ff <= -16'd4750;
        503: data_ff <= 16'd30638;
        504: data_ff <= 16'd7426;
        505: data_ff <= -16'd3046;
        506: data_ff <= 16'd1673;
        507: data_ff <= -16'd969;
        508: data_ff <= 16'd546;
        509: data_ff <= -16'd284;
        510: data_ff <= 16'd126;
        511: data_ff <= -16'd40;
        512: data_ff <= -16'd75;
        513: data_ff <= 16'd191;
        514: data_ff <= -16'd395;
        515: data_ff <= 16'd733;
        516: data_ff <= -16'd1296;
        517: data_ff <= 16'd2324;
        518: data_ff <= -16'd4855;
        519: data_ff <= 16'd30507;
        520: data_ff <= 16'd7689;
        521: data_ff <= -16'd3140;
        522: data_ff <= 16'd1723;
        523: data_ff <= -16'd997;
        524: data_ff <= 16'd562;
        525: data_ff <= -16'd292;
        526: data_ff <= 16'd130;
        527: data_ff <= -16'd41;
        528: data_ff <= -16'd77;
        529: data_ff <= 16'd196;
        530: data_ff <= -16'd404;
        531: data_ff <= 16'd751;
        532: data_ff <= -16'd1327;
        533: data_ff <= 16'd2378;
        534: data_ff <= -16'd4956;
        535: data_ff <= 16'd30372;
        536: data_ff <= 16'd7954;
        537: data_ff <= -16'd3234;
        538: data_ff <= 16'd1773;
        539: data_ff <= -16'd1026;
        540: data_ff <= 16'd578;
        541: data_ff <= -16'd300;
        542: data_ff <= 16'd134;
        543: data_ff <= -16'd43;
        544: data_ff <= -16'd79;
        545: data_ff <= 16'd200;
        546: data_ff <= -16'd414;
        547: data_ff <= 16'd768;
        548: data_ff <= -16'd1358;
        549: data_ff <= 16'd2431;
        550: data_ff <= -16'd5054;
        551: data_ff <= 16'd30233;
        552: data_ff <= 16'd8219;
        553: data_ff <= -16'd3328;
        554: data_ff <= 16'd1822;
        555: data_ff <= -16'd1054;
        556: data_ff <= 16'd594;
        557: data_ff <= -16'd309;
        558: data_ff <= 16'd138;
        559: data_ff <= -16'd44;
        560: data_ff <= -16'd80;
        561: data_ff <= 16'd204;
        562: data_ff <= -16'd423;
        563: data_ff <= 16'd785;
        564: data_ff <= -16'd1387;
        565: data_ff <= 16'd2482;
        566: data_ff <= -16'd5149;
        567: data_ff <= 16'd30091;
        568: data_ff <= 16'd8486;
        569: data_ff <= -16'd3421;
        570: data_ff <= 16'd1871;
        571: data_ff <= -16'd1081;
        572: data_ff <= 16'd610;
        573: data_ff <= -16'd317;
        574: data_ff <= 16'd141;
        575: data_ff <= -16'd46;
        576: data_ff <= -16'd82;
        577: data_ff <= 16'd208;
        578: data_ff <= -16'd432;
        579: data_ff <= 16'd802;
        580: data_ff <= -16'd1416;
        581: data_ff <= 16'd2532;
        582: data_ff <= -16'd5241;
        583: data_ff <= 16'd29945;
        584: data_ff <= 16'd8754;
        585: data_ff <= -16'd3513;
        586: data_ff <= 16'd1919;
        587: data_ff <= -16'd1109;
        588: data_ff <= 16'd625;
        589: data_ff <= -16'd325;
        590: data_ff <= 16'd145;
        591: data_ff <= -16'd47;
        592: data_ff <= -16'd83;
        593: data_ff <= 16'd213;
        594: data_ff <= -16'd440;
        595: data_ff <= 16'd818;
        596: data_ff <= -16'd1444;
        597: data_ff <= 16'd2580;
        598: data_ff <= -16'd5330;
        599: data_ff <= 16'd29795;
        600: data_ff <= 16'd9023;
        601: data_ff <= -16'd3605;
        602: data_ff <= 16'd1967;
        603: data_ff <= -16'd1136;
        604: data_ff <= 16'd641;
        605: data_ff <= -16'd333;
        606: data_ff <= 16'd149;
        607: data_ff <= -16'd48;
        608: data_ff <= -16'd85;
        609: data_ff <= 16'd216;
        610: data_ff <= -16'd449;
        611: data_ff <= 16'd834;
        612: data_ff <= -16'd1472;
        613: data_ff <= 16'd2627;
        614: data_ff <= -16'd5416;
        615: data_ff <= 16'd29642;
        616: data_ff <= 16'd9293;
        617: data_ff <= -16'd3696;
        618: data_ff <= 16'd2015;
        619: data_ff <= -16'd1164;
        620: data_ff <= 16'd656;
        621: data_ff <= -16'd342;
        622: data_ff <= 16'd153;
        623: data_ff <= -16'd50;
        624: data_ff <= -16'd86;
        625: data_ff <= 16'd220;
        626: data_ff <= -16'd457;
        627: data_ff <= 16'd849;
        628: data_ff <= -16'd1498;
        629: data_ff <= 16'd2673;
        630: data_ff <= -16'd5499;
        631: data_ff <= 16'd29485;
        632: data_ff <= 16'd9564;
        633: data_ff <= -16'd3787;
        634: data_ff <= 16'd2062;
        635: data_ff <= -16'd1190;
        636: data_ff <= 16'd671;
        637: data_ff <= -16'd350;
        638: data_ff <= 16'd157;
        639: data_ff <= -16'd51;
        640: data_ff <= -16'd87;
        641: data_ff <= 16'd224;
        642: data_ff <= -16'd465;
        643: data_ff <= 16'd864;
        644: data_ff <= -16'd1524;
        645: data_ff <= 16'd2717;
        646: data_ff <= -16'd5578;
        647: data_ff <= 16'd29325;
        648: data_ff <= 16'd9836;
        649: data_ff <= -16'd3877;
        650: data_ff <= 16'd2109;
        651: data_ff <= -16'd1217;
        652: data_ff <= 16'd686;
        653: data_ff <= -16'd358;
        654: data_ff <= 16'd160;
        655: data_ff <= -16'd52;
        656: data_ff <= -16'd89;
        657: data_ff <= 16'd227;
        658: data_ff <= -16'd472;
        659: data_ff <= 16'd878;
        660: data_ff <= -16'd1549;
        661: data_ff <= 16'd2760;
        662: data_ff <= -16'd5655;
        663: data_ff <= 16'd29162;
        664: data_ff <= 16'd10109;
        665: data_ff <= -16'd3966;
        666: data_ff <= 16'd2155;
        667: data_ff <= -16'd1243;
        668: data_ff <= 16'd701;
        669: data_ff <= -16'd365;
        670: data_ff <= 16'd164;
        671: data_ff <= -16'd54;
        672: data_ff <= -16'd90;
        673: data_ff <= 16'd231;
        674: data_ff <= -16'd479;
        675: data_ff <= 16'd892;
        676: data_ff <= -16'd1573;
        677: data_ff <= 16'd2802;
        678: data_ff <= -16'd5729;
        679: data_ff <= 16'd28994;
        680: data_ff <= 16'd10383;
        681: data_ff <= -16'd4054;
        682: data_ff <= 16'd2200;
        683: data_ff <= -16'd1269;
        684: data_ff <= 16'd716;
        685: data_ff <= -16'd373;
        686: data_ff <= 16'd168;
        687: data_ff <= -16'd55;
        688: data_ff <= -16'd91;
        689: data_ff <= 16'd234;
        690: data_ff <= -16'd487;
        691: data_ff <= 16'd905;
        692: data_ff <= -16'd1597;
        693: data_ff <= 16'd2842;
        694: data_ff <= -16'd5799;
        695: data_ff <= 16'd28824;
        696: data_ff <= 16'd10658;
        697: data_ff <= -16'd4142;
        698: data_ff <= 16'd2246;
        699: data_ff <= -16'd1295;
        700: data_ff <= 16'd730;
        701: data_ff <= -16'd381;
        702: data_ff <= 16'd172;
        703: data_ff <= -16'd57;
        704: data_ff <= -16'd92;
        705: data_ff <= 16'd237;
        706: data_ff <= -16'd493;
        707: data_ff <= 16'd918;
        708: data_ff <= -16'd1619;
        709: data_ff <= 16'd2880;
        710: data_ff <= -16'd5867;
        711: data_ff <= 16'd28650;
        712: data_ff <= 16'd10933;
        713: data_ff <= -16'd4229;
        714: data_ff <= 16'd2290;
        715: data_ff <= -16'd1320;
        716: data_ff <= 16'd745;
        717: data_ff <= -16'd389;
        718: data_ff <= 16'd175;
        719: data_ff <= -16'd58;
        720: data_ff <= -16'd93;
        721: data_ff <= 16'd240;
        722: data_ff <= -16'd500;
        723: data_ff <= 16'd930;
        724: data_ff <= -16'd1641;
        725: data_ff <= 16'd2918;
        726: data_ff <= -16'd5931;
        727: data_ff <= 16'd28473;
        728: data_ff <= 16'd11209;
        729: data_ff <= -16'd4314;
        730: data_ff <= 16'd2334;
        731: data_ff <= -16'd1345;
        732: data_ff <= 16'd759;
        733: data_ff <= -16'd396;
        734: data_ff <= 16'd179;
        735: data_ff <= -16'd59;
        736: data_ff <= -16'd94;
        737: data_ff <= 16'd243;
        738: data_ff <= -16'd506;
        739: data_ff <= 16'd942;
        740: data_ff <= -16'd1662;
        741: data_ff <= 16'd2953;
        742: data_ff <= -16'd5993;
        743: data_ff <= 16'd28293;
        744: data_ff <= 16'd11485;
        745: data_ff <= -16'd4399;
        746: data_ff <= 16'd2377;
        747: data_ff <= -16'd1370;
        748: data_ff <= 16'd773;
        749: data_ff <= -16'd404;
        750: data_ff <= 16'd182;
        751: data_ff <= -16'd61;
        752: data_ff <= -16'd95;
        753: data_ff <= 16'd246;
        754: data_ff <= -16'd512;
        755: data_ff <= 16'd954;
        756: data_ff <= -16'd1683;
        757: data_ff <= 16'd2988;
        758: data_ff <= -16'd6051;
        759: data_ff <= 16'd28109;
        760: data_ff <= 16'd11762;
        761: data_ff <= -16'd4483;
        762: data_ff <= 16'd2420;
        763: data_ff <= -16'd1394;
        764: data_ff <= 16'd786;
        765: data_ff <= -16'd411;
        766: data_ff <= 16'd186;
        767: data_ff <= -16'd62;
        768: data_ff <= -16'd96;
        769: data_ff <= 16'd248;
        770: data_ff <= -16'd518;
        771: data_ff <= 16'd965;
        772: data_ff <= -16'd1702;
        773: data_ff <= 16'd3021;
        774: data_ff <= -16'd6107;
        775: data_ff <= 16'd27922;
        776: data_ff <= 16'd12040;
        777: data_ff <= -16'd4566;
        778: data_ff <= 16'd2462;
        779: data_ff <= -16'd1418;
        780: data_ff <= 16'd800;
        781: data_ff <= -16'd418;
        782: data_ff <= 16'd189;
        783: data_ff <= -16'd63;
        784: data_ff <= -16'd96;
        785: data_ff <= 16'd251;
        786: data_ff <= -16'd524;
        787: data_ff <= 16'd976;
        788: data_ff <= -16'd1721;
        789: data_ff <= 16'd3052;
        790: data_ff <= -16'd6159;
        791: data_ff <= 16'd27732;
        792: data_ff <= 16'd12318;
        793: data_ff <= -16'd4648;
        794: data_ff <= 16'd2504;
        795: data_ff <= -16'd1441;
        796: data_ff <= 16'd813;
        797: data_ff <= -16'd425;
        798: data_ff <= 16'd193;
        799: data_ff <= -16'd65;
        800: data_ff <= -16'd97;
        801: data_ff <= 16'd253;
        802: data_ff <= -16'd529;
        803: data_ff <= 16'd986;
        804: data_ff <= -16'd1739;
        805: data_ff <= 16'd3082;
        806: data_ff <= -16'd6209;
        807: data_ff <= 16'd27539;
        808: data_ff <= 16'd12596;
        809: data_ff <= -16'd4728;
        810: data_ff <= 16'd2544;
        811: data_ff <= -16'd1464;
        812: data_ff <= 16'd826;
        813: data_ff <= -16'd433;
        814: data_ff <= 16'd196;
        815: data_ff <= -16'd66;
        816: data_ff <= -16'd98;
        817: data_ff <= 16'd255;
        818: data_ff <= -16'd534;
        819: data_ff <= 16'd996;
        820: data_ff <= -16'd1756;
        821: data_ff <= 16'd3111;
        822: data_ff <= -16'd6256;
        823: data_ff <= 16'd27343;
        824: data_ff <= 16'd12875;
        825: data_ff <= -16'd4808;
        826: data_ff <= 16'd2584;
        827: data_ff <= -16'd1487;
        828: data_ff <= 16'd839;
        829: data_ff <= -16'd439;
        830: data_ff <= 16'd199;
        831: data_ff <= -16'd67;
        832: data_ff <= -16'd99;
        833: data_ff <= 16'd258;
        834: data_ff <= -16'd539;
        835: data_ff <= 16'd1005;
        836: data_ff <= -16'd1772;
        837: data_ff <= 16'd3138;
        838: data_ff <= -16'd6299;
        839: data_ff <= 16'd27144;
        840: data_ff <= 16'd13154;
        841: data_ff <= -16'd4886;
        842: data_ff <= 16'd2623;
        843: data_ff <= -16'd1509;
        844: data_ff <= 16'd852;
        845: data_ff <= -16'd446;
        846: data_ff <= 16'd203;
        847: data_ff <= -16'd69;
        848: data_ff <= -16'd99;
        849: data_ff <= 16'd260;
        850: data_ff <= -16'd543;
        851: data_ff <= 16'd1014;
        852: data_ff <= -16'd1787;
        853: data_ff <= 16'd3164;
        854: data_ff <= -16'd6340;
        855: data_ff <= 16'd26942;
        856: data_ff <= 16'd13433;
        857: data_ff <= -16'd4963;
        858: data_ff <= 16'd2662;
        859: data_ff <= -16'd1531;
        860: data_ff <= 16'd864;
        861: data_ff <= -16'd453;
        862: data_ff <= 16'd206;
        863: data_ff <= -16'd70;
        864: data_ff <= -16'd100;
        865: data_ff <= 16'd261;
        866: data_ff <= -16'd548;
        867: data_ff <= 16'd1022;
        868: data_ff <= -16'd1802;
        869: data_ff <= 16'd3189;
        870: data_ff <= -16'd6378;
        871: data_ff <= 16'd26737;
        872: data_ff <= 16'd13712;
        873: data_ff <= -16'd5039;
        874: data_ff <= 16'd2700;
        875: data_ff <= -16'd1552;
        876: data_ff <= 16'd876;
        877: data_ff <= -16'd460;
        878: data_ff <= 16'd209;
        879: data_ff <= -16'd71;
        880: data_ff <= -16'd100;
        881: data_ff <= 16'd263;
        882: data_ff <= -16'd552;
        883: data_ff <= 16'd1030;
        884: data_ff <= -16'd1816;
        885: data_ff <= 16'd3211;
        886: data_ff <= -16'd6413;
        887: data_ff <= 16'd26530;
        888: data_ff <= 16'd13991;
        889: data_ff <= -16'd5114;
        890: data_ff <= 16'd2736;
        891: data_ff <= -16'd1573;
        892: data_ff <= 16'd888;
        893: data_ff <= -16'd466;
        894: data_ff <= 16'd212;
        895: data_ff <= -16'd72;
        896: data_ff <= -16'd101;
        897: data_ff <= 16'd265;
        898: data_ff <= -16'd555;
        899: data_ff <= 16'd1037;
        900: data_ff <= -16'd1829;
        901: data_ff <= 16'd3233;
        902: data_ff <= -16'd6445;
        903: data_ff <= 16'd26319;
        904: data_ff <= 16'd14271;
        905: data_ff <= -16'd5187;
        906: data_ff <= 16'd2773;
        907: data_ff <= -16'd1593;
        908: data_ff <= 16'd900;
        909: data_ff <= -16'd472;
        910: data_ff <= 16'd215;
        911: data_ff <= -16'd74;
        912: data_ff <= -16'd101;
        913: data_ff <= 16'd266;
        914: data_ff <= -16'd559;
        915: data_ff <= 16'd1044;
        916: data_ff <= -16'd1841;
        917: data_ff <= 16'd3253;
        918: data_ff <= -16'd6474;
        919: data_ff <= 16'd26106;
        920: data_ff <= 16'd14550;
        921: data_ff <= -16'd5259;
        922: data_ff <= 16'd2808;
        923: data_ff <= -16'd1613;
        924: data_ff <= 16'd911;
        925: data_ff <= -16'd478;
        926: data_ff <= 16'd218;
        927: data_ff <= -16'd75;
        928: data_ff <= -16'd101;
        929: data_ff <= 16'd267;
        930: data_ff <= -16'd562;
        931: data_ff <= 16'd1050;
        932: data_ff <= -16'd1852;
        933: data_ff <= 16'd3272;
        934: data_ff <= -16'd6501;
        935: data_ff <= 16'd25890;
        936: data_ff <= 16'd14829;
        937: data_ff <= -16'd5329;
        938: data_ff <= 16'd2842;
        939: data_ff <= -16'd1632;
        940: data_ff <= 16'd922;
        941: data_ff <= -16'd484;
        942: data_ff <= 16'd221;
        943: data_ff <= -16'd76;
        944: data_ff <= -16'd101;
        945: data_ff <= 16'd269;
        946: data_ff <= -16'd565;
        947: data_ff <= 16'd1056;
        948: data_ff <= -16'd1863;
        949: data_ff <= 16'd3289;
        950: data_ff <= -16'd6524;
        951: data_ff <= 16'd25671;
        952: data_ff <= 16'd15108;
        953: data_ff <= -16'd5398;
        954: data_ff <= 16'd2876;
        955: data_ff <= -16'd1651;
        956: data_ff <= 16'd933;
        957: data_ff <= -16'd490;
        958: data_ff <= 16'd224;
        959: data_ff <= -16'd77;
        960: data_ff <= -16'd102;
        961: data_ff <= 16'd270;
        962: data_ff <= -16'd568;
        963: data_ff <= 16'd1062;
        964: data_ff <= -16'd1873;
        965: data_ff <= 16'd3305;
        966: data_ff <= -16'd6545;
        967: data_ff <= 16'd25450;
        968: data_ff <= 16'd15387;
        969: data_ff <= -16'd5466;
        970: data_ff <= 16'd2908;
        971: data_ff <= -16'd1669;
        972: data_ff <= 16'd943;
        973: data_ff <= -16'd496;
        974: data_ff <= 16'd227;
        975: data_ff <= -16'd78;
        976: data_ff <= -16'd102;
        977: data_ff <= 16'd271;
        978: data_ff <= -16'd570;
        979: data_ff <= 16'd1067;
        980: data_ff <= -16'd1881;
        981: data_ff <= 16'd3319;
        982: data_ff <= -16'd6563;
        983: data_ff <= 16'd25226;
        984: data_ff <= 16'd15666;
        985: data_ff <= -16'd5532;
        986: data_ff <= 16'd2940;
        987: data_ff <= -16'd1687;
        988: data_ff <= 16'd953;
        989: data_ff <= -16'd502;
        990: data_ff <= 16'd230;
        991: data_ff <= -16'd80;
        992: data_ff <= -16'd102;
        993: data_ff <= 16'd272;
        994: data_ff <= -16'd573;
        995: data_ff <= 16'd1071;
        996: data_ff <= -16'd1890;
        997: data_ff <= 16'd3332;
        998: data_ff <= -16'd6578;
        999: data_ff <= 16'd25000;
        1000: data_ff <= 16'd15944;
        1001: data_ff <= -16'd5596;
        1002: data_ff <= 16'd2971;
        1003: data_ff <= -16'd1704;
        1004: data_ff <= 16'd963;
        1005: data_ff <= -16'd507;
        1006: data_ff <= 16'd233;
        1007: data_ff <= -16'd81;
        1008: data_ff <= -16'd102;
        1009: data_ff <= 16'd272;
        1010: data_ff <= -16'd575;
        1011: data_ff <= 16'd1076;
        1012: data_ff <= -16'd1897;
        1013: data_ff <= 16'd3344;
        1014: data_ff <= -16'd6591;
        1015: data_ff <= 16'd24771;
        1016: data_ff <= 16'd16222;
        1017: data_ff <= -16'd5659;
        1018: data_ff <= 16'd3001;
        1019: data_ff <= -16'd1721;
        1020: data_ff <= 16'd973;
        1021: data_ff <= -16'd512;
        1022: data_ff <= 16'd235;
        1023: data_ff <= -16'd82;
        1024: data_ff <= -16'd102;
        1025: data_ff <= 16'd273;
        1026: data_ff <= -16'd576;
        1027: data_ff <= 16'd1079;
        1028: data_ff <= -16'd1903;
        1029: data_ff <= 16'd3354;
        1030: data_ff <= -16'd6601;
        1031: data_ff <= 16'd24540;
        1032: data_ff <= 16'd16499;
        1033: data_ff <= -16'd5720;
        1034: data_ff <= 16'd3029;
        1035: data_ff <= -16'd1737;
        1036: data_ff <= 16'd982;
        1037: data_ff <= -16'd517;
        1038: data_ff <= 16'd238;
        1039: data_ff <= -16'd83;
        1040: data_ff <= -16'd102;
        1041: data_ff <= 16'd273;
        1042: data_ff <= -16'd578;
        1043: data_ff <= 16'd1082;
        1044: data_ff <= -16'd1909;
        1045: data_ff <= 16'd3363;
        1046: data_ff <= -16'd6608;
        1047: data_ff <= 16'd24307;
        1048: data_ff <= 16'd16776;
        1049: data_ff <= -16'd5779;
        1050: data_ff <= 16'd3057;
        1051: data_ff <= -16'd1752;
        1052: data_ff <= 16'd991;
        1053: data_ff <= -16'd522;
        1054: data_ff <= 16'd240;
        1055: data_ff <= -16'd84;
        1056: data_ff <= -16'd102;
        1057: data_ff <= 16'd274;
        1058: data_ff <= -16'd579;
        1059: data_ff <= 16'd1085;
        1060: data_ff <= -16'd1914;
        1061: data_ff <= 16'd3370;
        1062: data_ff <= -16'd6613;
        1063: data_ff <= 16'd24071;
        1064: data_ff <= 16'd17052;
        1065: data_ff <= -16'd5837;
        1066: data_ff <= 16'd3084;
        1067: data_ff <= -16'd1767;
        1068: data_ff <= 16'd999;
        1069: data_ff <= -16'd527;
        1070: data_ff <= 16'd243;
        1071: data_ff <= -16'd85;
        1072: data_ff <= -16'd102;
        1073: data_ff <= 16'd274;
        1074: data_ff <= -16'd580;
        1075: data_ff <= 16'd1087;
        1076: data_ff <= -16'd1918;
        1077: data_ff <= 16'd3376;
        1078: data_ff <= -16'd6615;
        1079: data_ff <= 16'd23833;
        1080: data_ff <= 16'd17328;
        1081: data_ff <= -16'd5893;
        1082: data_ff <= 16'd3110;
        1083: data_ff <= -16'd1781;
        1084: data_ff <= 16'd1007;
        1085: data_ff <= -16'd532;
        1086: data_ff <= 16'd245;
        1087: data_ff <= -16'd86;
        1088: data_ff <= -16'd102;
        1089: data_ff <= 16'd274;
        1090: data_ff <= -16'd581;
        1091: data_ff <= 16'd1089;
        1092: data_ff <= -16'd1922;
        1093: data_ff <= 16'd3381;
        1094: data_ff <= -16'd6614;
        1095: data_ff <= 16'd23593;
        1096: data_ff <= 16'd17603;
        1097: data_ff <= -16'd5947;
        1098: data_ff <= 16'd3135;
        1099: data_ff <= -16'd1795;
        1100: data_ff <= 16'd1015;
        1101: data_ff <= -16'd536;
        1102: data_ff <= 16'd247;
        1103: data_ff <= -16'd87;
        1104: data_ff <= -16'd101;
        1105: data_ff <= 16'd274;
        1106: data_ff <= -16'd581;
        1107: data_ff <= 16'd1091;
        1108: data_ff <= -16'd1924;
        1109: data_ff <= 16'd3384;
        1110: data_ff <= -16'd6611;
        1111: data_ff <= 16'd23351;
        1112: data_ff <= 16'd17877;
        1113: data_ff <= -16'd5999;
        1114: data_ff <= 16'd3158;
        1115: data_ff <= -16'd1808;
        1116: data_ff <= 16'd1023;
        1117: data_ff <= -16'd540;
        1118: data_ff <= 16'd250;
        1119: data_ff <= -16'd88;
        1120: data_ff <= -16'd101;
        1121: data_ff <= 16'd274;
        1122: data_ff <= -16'd582;
        1123: data_ff <= 16'd1092;
        1124: data_ff <= -16'd1926;
        1125: data_ff <= 16'd3386;
        1126: data_ff <= -16'd6605;
        1127: data_ff <= 16'd23106;
        1128: data_ff <= 16'd18150;
        1129: data_ff <= -16'd6050;
        1130: data_ff <= 16'd3181;
        1131: data_ff <= -16'd1821;
        1132: data_ff <= 16'd1030;
        1133: data_ff <= -16'd544;
        1134: data_ff <= 16'd252;
        1135: data_ff <= -16'd89;
        1136: data_ff <= -16'd101;
        1137: data_ff <= 16'd274;
        1138: data_ff <= -16'd582;
        1139: data_ff <= 16'd1092;
        1140: data_ff <= -16'd1927;
        1141: data_ff <= 16'd3387;
        1142: data_ff <= -16'd6597;
        1143: data_ff <= 16'd22860;
        1144: data_ff <= 16'd18422;
        1145: data_ff <= -16'd6098;
        1146: data_ff <= 16'd3203;
        1147: data_ff <= -16'd1832;
        1148: data_ff <= 16'd1037;
        1149: data_ff <= -16'd548;
        1150: data_ff <= 16'd254;
        1151: data_ff <= -16'd90;
        1152: data_ff <= -16'd101;
        1153: data_ff <= 16'd273;
        1154: data_ff <= -16'd581;
        1155: data_ff <= 16'd1092;
        1156: data_ff <= -16'd1927;
        1157: data_ff <= 16'd3386;
        1158: data_ff <= -16'd6586;
        1159: data_ff <= 16'd22612;
        1160: data_ff <= 16'd18694;
        1161: data_ff <= -16'd6145;
        1162: data_ff <= 16'd3223;
        1163: data_ff <= -16'd1843;
        1164: data_ff <= 16'd1043;
        1165: data_ff <= -16'd552;
        1166: data_ff <= 16'd256;
        1167: data_ff <= -16'd91;
        1168: data_ff <= -16'd100;
        1169: data_ff <= 16'd273;
        1170: data_ff <= -16'd581;
        1171: data_ff <= 16'd1092;
        1172: data_ff <= -16'd1927;
        1173: data_ff <= 16'd3384;
        1174: data_ff <= -16'd6572;
        1175: data_ff <= 16'd22362;
        1176: data_ff <= 16'd18964;
        1177: data_ff <= -16'd6189;
        1178: data_ff <= 16'd3242;
        1179: data_ff <= -16'd1854;
        1180: data_ff <= 16'd1049;
        1181: data_ff <= -16'd555;
        1182: data_ff <= 16'd258;
        1183: data_ff <= -16'd92;
        1184: data_ff <= -16'd100;
        1185: data_ff <= 16'd272;
        1186: data_ff <= -16'd580;
        1187: data_ff <= 16'd1091;
        1188: data_ff <= -16'd1926;
        1189: data_ff <= 16'd3381;
        1190: data_ff <= -16'd6557;
        1191: data_ff <= 16'd22110;
        1192: data_ff <= 16'd19234;
        1193: data_ff <= -16'd6232;
        1194: data_ff <= 16'd3260;
        1195: data_ff <= -16'd1864;
        1196: data_ff <= 16'd1055;
        1197: data_ff <= -16'd558;
        1198: data_ff <= 16'd259;
        1199: data_ff <= -16'd93;
        1200: data_ff <= -16'd99;
        1201: data_ff <= 16'd272;
        1202: data_ff <= -16'd579;
        1203: data_ff <= 16'd1090;
        1204: data_ff <= -16'd1924;
        1205: data_ff <= 16'd3376;
        1206: data_ff <= -16'd6539;
        1207: data_ff <= 16'd21856;
        1208: data_ff <= 16'd19502;
        1209: data_ff <= -16'd6272;
        1210: data_ff <= 16'd3277;
        1211: data_ff <= -16'd1873;
        1212: data_ff <= 16'd1060;
        1213: data_ff <= -16'd561;
        1214: data_ff <= 16'd261;
        1215: data_ff <= -16'd94;
        1216: data_ff <= -16'd99;
        1217: data_ff <= 16'd271;
        1218: data_ff <= -16'd578;
        1219: data_ff <= 16'd1088;
        1220: data_ff <= -16'd1921;
        1221: data_ff <= 16'd3370;
        1222: data_ff <= -16'd6518;
        1223: data_ff <= 16'd21601;
        1224: data_ff <= 16'd19769;
        1225: data_ff <= -16'd6311;
        1226: data_ff <= 16'd3293;
        1227: data_ff <= -16'd1881;
        1228: data_ff <= 16'd1065;
        1229: data_ff <= -16'd564;
        1230: data_ff <= 16'd263;
        1231: data_ff <= -16'd94;
        1232: data_ff <= -16'd98;
        1233: data_ff <= 16'd270;
        1234: data_ff <= -16'd577;
        1235: data_ff <= 16'd1086;
        1236: data_ff <= -16'd1917;
        1237: data_ff <= 16'd3363;
        1238: data_ff <= -16'd6495;
        1239: data_ff <= 16'd21343;
        1240: data_ff <= 16'd20035;
        1241: data_ff <= -16'd6347;
        1242: data_ff <= 16'd3308;
        1243: data_ff <= -16'd1889;
        1244: data_ff <= 16'd1069;
        1245: data_ff <= -16'd567;
        1246: data_ff <= 16'd264;
        1247: data_ff <= -16'd95;
        1248: data_ff <= -16'd98;
        1249: data_ff <= 16'd269;
        1250: data_ff <= -16'd575;
        1251: data_ff <= 16'd1084;
        1252: data_ff <= -16'd1913;
        1253: data_ff <= 16'd3354;
        1254: data_ff <= -16'd6470;
        1255: data_ff <= 16'd21085;
        1256: data_ff <= 16'd20300;
        1257: data_ff <= -16'd6381;
        1258: data_ff <= 16'd3321;
        1259: data_ff <= -16'd1896;
        1260: data_ff <= 16'd1074;
        1261: data_ff <= -16'd569;
        1262: data_ff <= 16'd265;
        1263: data_ff <= -16'd96;
        1264: data_ff <= -16'd97;
        1265: data_ff <= 16'd268;
        1266: data_ff <= -16'd574;
        1267: data_ff <= 16'd1081;
        1268: data_ff <= -16'd1908;
        1269: data_ff <= 16'd3345;
        1270: data_ff <= -16'd6443;
        1271: data_ff <= 16'd20824;
        1272: data_ff <= 16'd20563;
        1273: data_ff <= -16'd6413;
        1274: data_ff <= 16'd3334;
        1275: data_ff <= -16'd1903;
        1276: data_ff <= 16'd1077;
        1277: data_ff <= -16'd572;
        1278: data_ff <= 16'd267;
        1279: data_ff <= -16'd96;
        1280: data_ff <= -16'd96;
        1281: data_ff <= 16'd267;
        1282: data_ff <= -16'd572;
        1283: data_ff <= 16'd1077;
        1284: data_ff <= -16'd1903;
        1285: data_ff <= 16'd3334;
        1286: data_ff <= -16'd6413;
        1287: data_ff <= 16'd20563;
        1288: data_ff <= 16'd20824;
        1289: data_ff <= -16'd6443;
        1290: data_ff <= 16'd3345;
        1291: data_ff <= -16'd1908;
        1292: data_ff <= 16'd1081;
        1293: data_ff <= -16'd574;
        1294: data_ff <= 16'd268;
        1295: data_ff <= -16'd97;
        1296: data_ff <= -16'd96;
        1297: data_ff <= 16'd265;
        1298: data_ff <= -16'd569;
        1299: data_ff <= 16'd1074;
        1300: data_ff <= -16'd1896;
        1301: data_ff <= 16'd3321;
        1302: data_ff <= -16'd6381;
        1303: data_ff <= 16'd20300;
        1304: data_ff <= 16'd21085;
        1305: data_ff <= -16'd6470;
        1306: data_ff <= 16'd3354;
        1307: data_ff <= -16'd1913;
        1308: data_ff <= 16'd1084;
        1309: data_ff <= -16'd575;
        1310: data_ff <= 16'd269;
        1311: data_ff <= -16'd98;
        1312: data_ff <= -16'd95;
        1313: data_ff <= 16'd264;
        1314: data_ff <= -16'd567;
        1315: data_ff <= 16'd1069;
        1316: data_ff <= -16'd1889;
        1317: data_ff <= 16'd3308;
        1318: data_ff <= -16'd6347;
        1319: data_ff <= 16'd20035;
        1320: data_ff <= 16'd21343;
        1321: data_ff <= -16'd6495;
        1322: data_ff <= 16'd3363;
        1323: data_ff <= -16'd1917;
        1324: data_ff <= 16'd1086;
        1325: data_ff <= -16'd577;
        1326: data_ff <= 16'd270;
        1327: data_ff <= -16'd98;
        1328: data_ff <= -16'd94;
        1329: data_ff <= 16'd263;
        1330: data_ff <= -16'd564;
        1331: data_ff <= 16'd1065;
        1332: data_ff <= -16'd1881;
        1333: data_ff <= 16'd3293;
        1334: data_ff <= -16'd6311;
        1335: data_ff <= 16'd19769;
        1336: data_ff <= 16'd21601;
        1337: data_ff <= -16'd6518;
        1338: data_ff <= 16'd3370;
        1339: data_ff <= -16'd1921;
        1340: data_ff <= 16'd1088;
        1341: data_ff <= -16'd578;
        1342: data_ff <= 16'd271;
        1343: data_ff <= -16'd99;
        1344: data_ff <= -16'd94;
        1345: data_ff <= 16'd261;
        1346: data_ff <= -16'd561;
        1347: data_ff <= 16'd1060;
        1348: data_ff <= -16'd1873;
        1349: data_ff <= 16'd3277;
        1350: data_ff <= -16'd6272;
        1351: data_ff <= 16'd19502;
        1352: data_ff <= 16'd21856;
        1353: data_ff <= -16'd6539;
        1354: data_ff <= 16'd3376;
        1355: data_ff <= -16'd1924;
        1356: data_ff <= 16'd1090;
        1357: data_ff <= -16'd579;
        1358: data_ff <= 16'd272;
        1359: data_ff <= -16'd99;
        1360: data_ff <= -16'd93;
        1361: data_ff <= 16'd259;
        1362: data_ff <= -16'd558;
        1363: data_ff <= 16'd1055;
        1364: data_ff <= -16'd1864;
        1365: data_ff <= 16'd3260;
        1366: data_ff <= -16'd6232;
        1367: data_ff <= 16'd19234;
        1368: data_ff <= 16'd22110;
        1369: data_ff <= -16'd6557;
        1370: data_ff <= 16'd3381;
        1371: data_ff <= -16'd1926;
        1372: data_ff <= 16'd1091;
        1373: data_ff <= -16'd580;
        1374: data_ff <= 16'd272;
        1375: data_ff <= -16'd100;
        1376: data_ff <= -16'd92;
        1377: data_ff <= 16'd258;
        1378: data_ff <= -16'd555;
        1379: data_ff <= 16'd1049;
        1380: data_ff <= -16'd1854;
        1381: data_ff <= 16'd3242;
        1382: data_ff <= -16'd6189;
        1383: data_ff <= 16'd18964;
        1384: data_ff <= 16'd22362;
        1385: data_ff <= -16'd6572;
        1386: data_ff <= 16'd3384;
        1387: data_ff <= -16'd1927;
        1388: data_ff <= 16'd1092;
        1389: data_ff <= -16'd581;
        1390: data_ff <= 16'd273;
        1391: data_ff <= -16'd100;
        1392: data_ff <= -16'd91;
        1393: data_ff <= 16'd256;
        1394: data_ff <= -16'd552;
        1395: data_ff <= 16'd1043;
        1396: data_ff <= -16'd1843;
        1397: data_ff <= 16'd3223;
        1398: data_ff <= -16'd6145;
        1399: data_ff <= 16'd18694;
        1400: data_ff <= 16'd22612;
        1401: data_ff <= -16'd6586;
        1402: data_ff <= 16'd3386;
        1403: data_ff <= -16'd1927;
        1404: data_ff <= 16'd1092;
        1405: data_ff <= -16'd581;
        1406: data_ff <= 16'd273;
        1407: data_ff <= -16'd101;
        1408: data_ff <= -16'd90;
        1409: data_ff <= 16'd254;
        1410: data_ff <= -16'd548;
        1411: data_ff <= 16'd1037;
        1412: data_ff <= -16'd1832;
        1413: data_ff <= 16'd3203;
        1414: data_ff <= -16'd6098;
        1415: data_ff <= 16'd18422;
        1416: data_ff <= 16'd22860;
        1417: data_ff <= -16'd6597;
        1418: data_ff <= 16'd3387;
        1419: data_ff <= -16'd1927;
        1420: data_ff <= 16'd1092;
        1421: data_ff <= -16'd582;
        1422: data_ff <= 16'd274;
        1423: data_ff <= -16'd101;
        1424: data_ff <= -16'd89;
        1425: data_ff <= 16'd252;
        1426: data_ff <= -16'd544;
        1427: data_ff <= 16'd1030;
        1428: data_ff <= -16'd1821;
        1429: data_ff <= 16'd3181;
        1430: data_ff <= -16'd6050;
        1431: data_ff <= 16'd18150;
        1432: data_ff <= 16'd23106;
        1433: data_ff <= -16'd6605;
        1434: data_ff <= 16'd3386;
        1435: data_ff <= -16'd1926;
        1436: data_ff <= 16'd1092;
        1437: data_ff <= -16'd582;
        1438: data_ff <= 16'd274;
        1439: data_ff <= -16'd101;
        1440: data_ff <= -16'd88;
        1441: data_ff <= 16'd250;
        1442: data_ff <= -16'd540;
        1443: data_ff <= 16'd1023;
        1444: data_ff <= -16'd1808;
        1445: data_ff <= 16'd3158;
        1446: data_ff <= -16'd5999;
        1447: data_ff <= 16'd17877;
        1448: data_ff <= 16'd23351;
        1449: data_ff <= -16'd6611;
        1450: data_ff <= 16'd3384;
        1451: data_ff <= -16'd1924;
        1452: data_ff <= 16'd1091;
        1453: data_ff <= -16'd581;
        1454: data_ff <= 16'd274;
        1455: data_ff <= -16'd101;
        1456: data_ff <= -16'd87;
        1457: data_ff <= 16'd247;
        1458: data_ff <= -16'd536;
        1459: data_ff <= 16'd1015;
        1460: data_ff <= -16'd1795;
        1461: data_ff <= 16'd3135;
        1462: data_ff <= -16'd5947;
        1463: data_ff <= 16'd17603;
        1464: data_ff <= 16'd23593;
        1465: data_ff <= -16'd6614;
        1466: data_ff <= 16'd3381;
        1467: data_ff <= -16'd1922;
        1468: data_ff <= 16'd1089;
        1469: data_ff <= -16'd581;
        1470: data_ff <= 16'd274;
        1471: data_ff <= -16'd102;
        1472: data_ff <= -16'd86;
        1473: data_ff <= 16'd245;
        1474: data_ff <= -16'd532;
        1475: data_ff <= 16'd1007;
        1476: data_ff <= -16'd1781;
        1477: data_ff <= 16'd3110;
        1478: data_ff <= -16'd5893;
        1479: data_ff <= 16'd17328;
        1480: data_ff <= 16'd23833;
        1481: data_ff <= -16'd6615;
        1482: data_ff <= 16'd3376;
        1483: data_ff <= -16'd1918;
        1484: data_ff <= 16'd1087;
        1485: data_ff <= -16'd580;
        1486: data_ff <= 16'd274;
        1487: data_ff <= -16'd102;
        1488: data_ff <= -16'd85;
        1489: data_ff <= 16'd243;
        1490: data_ff <= -16'd527;
        1491: data_ff <= 16'd999;
        1492: data_ff <= -16'd1767;
        1493: data_ff <= 16'd3084;
        1494: data_ff <= -16'd5837;
        1495: data_ff <= 16'd17052;
        1496: data_ff <= 16'd24071;
        1497: data_ff <= -16'd6613;
        1498: data_ff <= 16'd3370;
        1499: data_ff <= -16'd1914;
        1500: data_ff <= 16'd1085;
        1501: data_ff <= -16'd579;
        1502: data_ff <= 16'd274;
        1503: data_ff <= -16'd102;
        1504: data_ff <= -16'd84;
        1505: data_ff <= 16'd240;
        1506: data_ff <= -16'd522;
        1507: data_ff <= 16'd991;
        1508: data_ff <= -16'd1752;
        1509: data_ff <= 16'd3057;
        1510: data_ff <= -16'd5779;
        1511: data_ff <= 16'd16776;
        1512: data_ff <= 16'd24307;
        1513: data_ff <= -16'd6608;
        1514: data_ff <= 16'd3363;
        1515: data_ff <= -16'd1909;
        1516: data_ff <= 16'd1082;
        1517: data_ff <= -16'd578;
        1518: data_ff <= 16'd273;
        1519: data_ff <= -16'd102;
        1520: data_ff <= -16'd83;
        1521: data_ff <= 16'd238;
        1522: data_ff <= -16'd517;
        1523: data_ff <= 16'd982;
        1524: data_ff <= -16'd1737;
        1525: data_ff <= 16'd3029;
        1526: data_ff <= -16'd5720;
        1527: data_ff <= 16'd16499;
        1528: data_ff <= 16'd24540;
        1529: data_ff <= -16'd6601;
        1530: data_ff <= 16'd3354;
        1531: data_ff <= -16'd1903;
        1532: data_ff <= 16'd1079;
        1533: data_ff <= -16'd576;
        1534: data_ff <= 16'd273;
        1535: data_ff <= -16'd102;
        1536: data_ff <= -16'd82;
        1537: data_ff <= 16'd235;
        1538: data_ff <= -16'd512;
        1539: data_ff <= 16'd973;
        1540: data_ff <= -16'd1721;
        1541: data_ff <= 16'd3001;
        1542: data_ff <= -16'd5659;
        1543: data_ff <= 16'd16222;
        1544: data_ff <= 16'd24771;
        1545: data_ff <= -16'd6591;
        1546: data_ff <= 16'd3344;
        1547: data_ff <= -16'd1897;
        1548: data_ff <= 16'd1076;
        1549: data_ff <= -16'd575;
        1550: data_ff <= 16'd272;
        1551: data_ff <= -16'd102;
        1552: data_ff <= -16'd81;
        1553: data_ff <= 16'd233;
        1554: data_ff <= -16'd507;
        1555: data_ff <= 16'd963;
        1556: data_ff <= -16'd1704;
        1557: data_ff <= 16'd2971;
        1558: data_ff <= -16'd5596;
        1559: data_ff <= 16'd15944;
        1560: data_ff <= 16'd25000;
        1561: data_ff <= -16'd6578;
        1562: data_ff <= 16'd3332;
        1563: data_ff <= -16'd1890;
        1564: data_ff <= 16'd1071;
        1565: data_ff <= -16'd573;
        1566: data_ff <= 16'd272;
        1567: data_ff <= -16'd102;
        1568: data_ff <= -16'd80;
        1569: data_ff <= 16'd230;
        1570: data_ff <= -16'd502;
        1571: data_ff <= 16'd953;
        1572: data_ff <= -16'd1687;
        1573: data_ff <= 16'd2940;
        1574: data_ff <= -16'd5532;
        1575: data_ff <= 16'd15666;
        1576: data_ff <= 16'd25226;
        1577: data_ff <= -16'd6563;
        1578: data_ff <= 16'd3319;
        1579: data_ff <= -16'd1881;
        1580: data_ff <= 16'd1067;
        1581: data_ff <= -16'd570;
        1582: data_ff <= 16'd271;
        1583: data_ff <= -16'd102;
        1584: data_ff <= -16'd78;
        1585: data_ff <= 16'd227;
        1586: data_ff <= -16'd496;
        1587: data_ff <= 16'd943;
        1588: data_ff <= -16'd1669;
        1589: data_ff <= 16'd2908;
        1590: data_ff <= -16'd5466;
        1591: data_ff <= 16'd15387;
        1592: data_ff <= 16'd25450;
        1593: data_ff <= -16'd6545;
        1594: data_ff <= 16'd3305;
        1595: data_ff <= -16'd1873;
        1596: data_ff <= 16'd1062;
        1597: data_ff <= -16'd568;
        1598: data_ff <= 16'd270;
        1599: data_ff <= -16'd102;
        1600: data_ff <= -16'd77;
        1601: data_ff <= 16'd224;
        1602: data_ff <= -16'd490;
        1603: data_ff <= 16'd933;
        1604: data_ff <= -16'd1651;
        1605: data_ff <= 16'd2876;
        1606: data_ff <= -16'd5398;
        1607: data_ff <= 16'd15108;
        1608: data_ff <= 16'd25671;
        1609: data_ff <= -16'd6524;
        1610: data_ff <= 16'd3289;
        1611: data_ff <= -16'd1863;
        1612: data_ff <= 16'd1056;
        1613: data_ff <= -16'd565;
        1614: data_ff <= 16'd269;
        1615: data_ff <= -16'd101;
        1616: data_ff <= -16'd76;
        1617: data_ff <= 16'd221;
        1618: data_ff <= -16'd484;
        1619: data_ff <= 16'd922;
        1620: data_ff <= -16'd1632;
        1621: data_ff <= 16'd2842;
        1622: data_ff <= -16'd5329;
        1623: data_ff <= 16'd14829;
        1624: data_ff <= 16'd25890;
        1625: data_ff <= -16'd6501;
        1626: data_ff <= 16'd3272;
        1627: data_ff <= -16'd1852;
        1628: data_ff <= 16'd1050;
        1629: data_ff <= -16'd562;
        1630: data_ff <= 16'd267;
        1631: data_ff <= -16'd101;
        1632: data_ff <= -16'd75;
        1633: data_ff <= 16'd218;
        1634: data_ff <= -16'd478;
        1635: data_ff <= 16'd911;
        1636: data_ff <= -16'd1613;
        1637: data_ff <= 16'd2808;
        1638: data_ff <= -16'd5259;
        1639: data_ff <= 16'd14550;
        1640: data_ff <= 16'd26106;
        1641: data_ff <= -16'd6474;
        1642: data_ff <= 16'd3253;
        1643: data_ff <= -16'd1841;
        1644: data_ff <= 16'd1044;
        1645: data_ff <= -16'd559;
        1646: data_ff <= 16'd266;
        1647: data_ff <= -16'd101;
        1648: data_ff <= -16'd74;
        1649: data_ff <= 16'd215;
        1650: data_ff <= -16'd472;
        1651: data_ff <= 16'd900;
        1652: data_ff <= -16'd1593;
        1653: data_ff <= 16'd2773;
        1654: data_ff <= -16'd5187;
        1655: data_ff <= 16'd14271;
        1656: data_ff <= 16'd26319;
        1657: data_ff <= -16'd6445;
        1658: data_ff <= 16'd3233;
        1659: data_ff <= -16'd1829;
        1660: data_ff <= 16'd1037;
        1661: data_ff <= -16'd555;
        1662: data_ff <= 16'd265;
        1663: data_ff <= -16'd101;
        1664: data_ff <= -16'd72;
        1665: data_ff <= 16'd212;
        1666: data_ff <= -16'd466;
        1667: data_ff <= 16'd888;
        1668: data_ff <= -16'd1573;
        1669: data_ff <= 16'd2736;
        1670: data_ff <= -16'd5114;
        1671: data_ff <= 16'd13991;
        1672: data_ff <= 16'd26530;
        1673: data_ff <= -16'd6413;
        1674: data_ff <= 16'd3211;
        1675: data_ff <= -16'd1816;
        1676: data_ff <= 16'd1030;
        1677: data_ff <= -16'd552;
        1678: data_ff <= 16'd263;
        1679: data_ff <= -16'd100;
        1680: data_ff <= -16'd71;
        1681: data_ff <= 16'd209;
        1682: data_ff <= -16'd460;
        1683: data_ff <= 16'd876;
        1684: data_ff <= -16'd1552;
        1685: data_ff <= 16'd2700;
        1686: data_ff <= -16'd5039;
        1687: data_ff <= 16'd13712;
        1688: data_ff <= 16'd26737;
        1689: data_ff <= -16'd6378;
        1690: data_ff <= 16'd3189;
        1691: data_ff <= -16'd1802;
        1692: data_ff <= 16'd1022;
        1693: data_ff <= -16'd548;
        1694: data_ff <= 16'd261;
        1695: data_ff <= -16'd100;
        1696: data_ff <= -16'd70;
        1697: data_ff <= 16'd206;
        1698: data_ff <= -16'd453;
        1699: data_ff <= 16'd864;
        1700: data_ff <= -16'd1531;
        1701: data_ff <= 16'd2662;
        1702: data_ff <= -16'd4963;
        1703: data_ff <= 16'd13433;
        1704: data_ff <= 16'd26942;
        1705: data_ff <= -16'd6340;
        1706: data_ff <= 16'd3164;
        1707: data_ff <= -16'd1787;
        1708: data_ff <= 16'd1014;
        1709: data_ff <= -16'd543;
        1710: data_ff <= 16'd260;
        1711: data_ff <= -16'd99;
        1712: data_ff <= -16'd69;
        1713: data_ff <= 16'd203;
        1714: data_ff <= -16'd446;
        1715: data_ff <= 16'd852;
        1716: data_ff <= -16'd1509;
        1717: data_ff <= 16'd2623;
        1718: data_ff <= -16'd4886;
        1719: data_ff <= 16'd13154;
        1720: data_ff <= 16'd27144;
        1721: data_ff <= -16'd6299;
        1722: data_ff <= 16'd3138;
        1723: data_ff <= -16'd1772;
        1724: data_ff <= 16'd1005;
        1725: data_ff <= -16'd539;
        1726: data_ff <= 16'd258;
        1727: data_ff <= -16'd99;
        1728: data_ff <= -16'd67;
        1729: data_ff <= 16'd199;
        1730: data_ff <= -16'd439;
        1731: data_ff <= 16'd839;
        1732: data_ff <= -16'd1487;
        1733: data_ff <= 16'd2584;
        1734: data_ff <= -16'd4808;
        1735: data_ff <= 16'd12875;
        1736: data_ff <= 16'd27343;
        1737: data_ff <= -16'd6256;
        1738: data_ff <= 16'd3111;
        1739: data_ff <= -16'd1756;
        1740: data_ff <= 16'd996;
        1741: data_ff <= -16'd534;
        1742: data_ff <= 16'd255;
        1743: data_ff <= -16'd98;
        1744: data_ff <= -16'd66;
        1745: data_ff <= 16'd196;
        1746: data_ff <= -16'd433;
        1747: data_ff <= 16'd826;
        1748: data_ff <= -16'd1464;
        1749: data_ff <= 16'd2544;
        1750: data_ff <= -16'd4728;
        1751: data_ff <= 16'd12596;
        1752: data_ff <= 16'd27539;
        1753: data_ff <= -16'd6209;
        1754: data_ff <= 16'd3082;
        1755: data_ff <= -16'd1739;
        1756: data_ff <= 16'd986;
        1757: data_ff <= -16'd529;
        1758: data_ff <= 16'd253;
        1759: data_ff <= -16'd97;
        1760: data_ff <= -16'd65;
        1761: data_ff <= 16'd193;
        1762: data_ff <= -16'd425;
        1763: data_ff <= 16'd813;
        1764: data_ff <= -16'd1441;
        1765: data_ff <= 16'd2504;
        1766: data_ff <= -16'd4648;
        1767: data_ff <= 16'd12318;
        1768: data_ff <= 16'd27732;
        1769: data_ff <= -16'd6159;
        1770: data_ff <= 16'd3052;
        1771: data_ff <= -16'd1721;
        1772: data_ff <= 16'd976;
        1773: data_ff <= -16'd524;
        1774: data_ff <= 16'd251;
        1775: data_ff <= -16'd96;
        1776: data_ff <= -16'd63;
        1777: data_ff <= 16'd189;
        1778: data_ff <= -16'd418;
        1779: data_ff <= 16'd800;
        1780: data_ff <= -16'd1418;
        1781: data_ff <= 16'd2462;
        1782: data_ff <= -16'd4566;
        1783: data_ff <= 16'd12040;
        1784: data_ff <= 16'd27922;
        1785: data_ff <= -16'd6107;
        1786: data_ff <= 16'd3021;
        1787: data_ff <= -16'd1702;
        1788: data_ff <= 16'd965;
        1789: data_ff <= -16'd518;
        1790: data_ff <= 16'd248;
        1791: data_ff <= -16'd96;
        1792: data_ff <= -16'd62;
        1793: data_ff <= 16'd186;
        1794: data_ff <= -16'd411;
        1795: data_ff <= 16'd786;
        1796: data_ff <= -16'd1394;
        1797: data_ff <= 16'd2420;
        1798: data_ff <= -16'd4483;
        1799: data_ff <= 16'd11762;
        1800: data_ff <= 16'd28109;
        1801: data_ff <= -16'd6051;
        1802: data_ff <= 16'd2988;
        1803: data_ff <= -16'd1683;
        1804: data_ff <= 16'd954;
        1805: data_ff <= -16'd512;
        1806: data_ff <= 16'd246;
        1807: data_ff <= -16'd95;
        1808: data_ff <= -16'd61;
        1809: data_ff <= 16'd182;
        1810: data_ff <= -16'd404;
        1811: data_ff <= 16'd773;
        1812: data_ff <= -16'd1370;
        1813: data_ff <= 16'd2377;
        1814: data_ff <= -16'd4399;
        1815: data_ff <= 16'd11485;
        1816: data_ff <= 16'd28293;
        1817: data_ff <= -16'd5993;
        1818: data_ff <= 16'd2953;
        1819: data_ff <= -16'd1662;
        1820: data_ff <= 16'd942;
        1821: data_ff <= -16'd506;
        1822: data_ff <= 16'd243;
        1823: data_ff <= -16'd94;
        1824: data_ff <= -16'd59;
        1825: data_ff <= 16'd179;
        1826: data_ff <= -16'd396;
        1827: data_ff <= 16'd759;
        1828: data_ff <= -16'd1345;
        1829: data_ff <= 16'd2334;
        1830: data_ff <= -16'd4314;
        1831: data_ff <= 16'd11209;
        1832: data_ff <= 16'd28473;
        1833: data_ff <= -16'd5931;
        1834: data_ff <= 16'd2918;
        1835: data_ff <= -16'd1641;
        1836: data_ff <= 16'd930;
        1837: data_ff <= -16'd500;
        1838: data_ff <= 16'd240;
        1839: data_ff <= -16'd93;
        1840: data_ff <= -16'd58;
        1841: data_ff <= 16'd175;
        1842: data_ff <= -16'd389;
        1843: data_ff <= 16'd745;
        1844: data_ff <= -16'd1320;
        1845: data_ff <= 16'd2290;
        1846: data_ff <= -16'd4229;
        1847: data_ff <= 16'd10933;
        1848: data_ff <= 16'd28650;
        1849: data_ff <= -16'd5867;
        1850: data_ff <= 16'd2880;
        1851: data_ff <= -16'd1619;
        1852: data_ff <= 16'd918;
        1853: data_ff <= -16'd493;
        1854: data_ff <= 16'd237;
        1855: data_ff <= -16'd92;
        1856: data_ff <= -16'd57;
        1857: data_ff <= 16'd172;
        1858: data_ff <= -16'd381;
        1859: data_ff <= 16'd730;
        1860: data_ff <= -16'd1295;
        1861: data_ff <= 16'd2246;
        1862: data_ff <= -16'd4142;
        1863: data_ff <= 16'd10658;
        1864: data_ff <= 16'd28824;
        1865: data_ff <= -16'd5799;
        1866: data_ff <= 16'd2842;
        1867: data_ff <= -16'd1597;
        1868: data_ff <= 16'd905;
        1869: data_ff <= -16'd487;
        1870: data_ff <= 16'd234;
        1871: data_ff <= -16'd91;
        1872: data_ff <= -16'd55;
        1873: data_ff <= 16'd168;
        1874: data_ff <= -16'd373;
        1875: data_ff <= 16'd716;
        1876: data_ff <= -16'd1269;
        1877: data_ff <= 16'd2200;
        1878: data_ff <= -16'd4054;
        1879: data_ff <= 16'd10383;
        1880: data_ff <= 16'd28994;
        1881: data_ff <= -16'd5729;
        1882: data_ff <= 16'd2802;
        1883: data_ff <= -16'd1573;
        1884: data_ff <= 16'd892;
        1885: data_ff <= -16'd479;
        1886: data_ff <= 16'd231;
        1887: data_ff <= -16'd90;
        1888: data_ff <= -16'd54;
        1889: data_ff <= 16'd164;
        1890: data_ff <= -16'd365;
        1891: data_ff <= 16'd701;
        1892: data_ff <= -16'd1243;
        1893: data_ff <= 16'd2155;
        1894: data_ff <= -16'd3966;
        1895: data_ff <= 16'd10109;
        1896: data_ff <= 16'd29162;
        1897: data_ff <= -16'd5655;
        1898: data_ff <= 16'd2760;
        1899: data_ff <= -16'd1549;
        1900: data_ff <= 16'd878;
        1901: data_ff <= -16'd472;
        1902: data_ff <= 16'd227;
        1903: data_ff <= -16'd89;
        1904: data_ff <= -16'd52;
        1905: data_ff <= 16'd160;
        1906: data_ff <= -16'd358;
        1907: data_ff <= 16'd686;
        1908: data_ff <= -16'd1217;
        1909: data_ff <= 16'd2109;
        1910: data_ff <= -16'd3877;
        1911: data_ff <= 16'd9836;
        1912: data_ff <= 16'd29325;
        1913: data_ff <= -16'd5578;
        1914: data_ff <= 16'd2717;
        1915: data_ff <= -16'd1524;
        1916: data_ff <= 16'd864;
        1917: data_ff <= -16'd465;
        1918: data_ff <= 16'd224;
        1919: data_ff <= -16'd87;
        1920: data_ff <= -16'd51;
        1921: data_ff <= 16'd157;
        1922: data_ff <= -16'd350;
        1923: data_ff <= 16'd671;
        1924: data_ff <= -16'd1190;
        1925: data_ff <= 16'd2062;
        1926: data_ff <= -16'd3787;
        1927: data_ff <= 16'd9564;
        1928: data_ff <= 16'd29485;
        1929: data_ff <= -16'd5499;
        1930: data_ff <= 16'd2673;
        1931: data_ff <= -16'd1498;
        1932: data_ff <= 16'd849;
        1933: data_ff <= -16'd457;
        1934: data_ff <= 16'd220;
        1935: data_ff <= -16'd86;
        1936: data_ff <= -16'd50;
        1937: data_ff <= 16'd153;
        1938: data_ff <= -16'd342;
        1939: data_ff <= 16'd656;
        1940: data_ff <= -16'd1164;
        1941: data_ff <= 16'd2015;
        1942: data_ff <= -16'd3696;
        1943: data_ff <= 16'd9293;
        1944: data_ff <= 16'd29642;
        1945: data_ff <= -16'd5416;
        1946: data_ff <= 16'd2627;
        1947: data_ff <= -16'd1472;
        1948: data_ff <= 16'd834;
        1949: data_ff <= -16'd449;
        1950: data_ff <= 16'd216;
        1951: data_ff <= -16'd85;
        1952: data_ff <= -16'd48;
        1953: data_ff <= 16'd149;
        1954: data_ff <= -16'd333;
        1955: data_ff <= 16'd641;
        1956: data_ff <= -16'd1136;
        1957: data_ff <= 16'd1967;
        1958: data_ff <= -16'd3605;
        1959: data_ff <= 16'd9023;
        1960: data_ff <= 16'd29795;
        1961: data_ff <= -16'd5330;
        1962: data_ff <= 16'd2580;
        1963: data_ff <= -16'd1444;
        1964: data_ff <= 16'd818;
        1965: data_ff <= -16'd440;
        1966: data_ff <= 16'd213;
        1967: data_ff <= -16'd83;
        1968: data_ff <= -16'd47;
        1969: data_ff <= 16'd145;
        1970: data_ff <= -16'd325;
        1971: data_ff <= 16'd625;
        1972: data_ff <= -16'd1109;
        1973: data_ff <= 16'd1919;
        1974: data_ff <= -16'd3513;
        1975: data_ff <= 16'd8754;
        1976: data_ff <= 16'd29945;
        1977: data_ff <= -16'd5241;
        1978: data_ff <= 16'd2532;
        1979: data_ff <= -16'd1416;
        1980: data_ff <= 16'd802;
        1981: data_ff <= -16'd432;
        1982: data_ff <= 16'd208;
        1983: data_ff <= -16'd82;
        1984: data_ff <= -16'd46;
        1985: data_ff <= 16'd141;
        1986: data_ff <= -16'd317;
        1987: data_ff <= 16'd610;
        1988: data_ff <= -16'd1081;
        1989: data_ff <= 16'd1871;
        1990: data_ff <= -16'd3421;
        1991: data_ff <= 16'd8486;
        1992: data_ff <= 16'd30091;
        1993: data_ff <= -16'd5149;
        1994: data_ff <= 16'd2482;
        1995: data_ff <= -16'd1387;
        1996: data_ff <= 16'd785;
        1997: data_ff <= -16'd423;
        1998: data_ff <= 16'd204;
        1999: data_ff <= -16'd80;
        2000: data_ff <= -16'd44;
        2001: data_ff <= 16'd138;
        2002: data_ff <= -16'd309;
        2003: data_ff <= 16'd594;
        2004: data_ff <= -16'd1054;
        2005: data_ff <= 16'd1822;
        2006: data_ff <= -16'd3328;
        2007: data_ff <= 16'd8219;
        2008: data_ff <= 16'd30233;
        2009: data_ff <= -16'd5054;
        2010: data_ff <= 16'd2431;
        2011: data_ff <= -16'd1358;
        2012: data_ff <= 16'd768;
        2013: data_ff <= -16'd414;
        2014: data_ff <= 16'd200;
        2015: data_ff <= -16'd79;
        2016: data_ff <= -16'd43;
        2017: data_ff <= 16'd134;
        2018: data_ff <= -16'd300;
        2019: data_ff <= 16'd578;
        2020: data_ff <= -16'd1026;
        2021: data_ff <= 16'd1773;
        2022: data_ff <= -16'd3234;
        2023: data_ff <= 16'd7954;
        2024: data_ff <= 16'd30372;
        2025: data_ff <= -16'd4956;
        2026: data_ff <= 16'd2378;
        2027: data_ff <= -16'd1327;
        2028: data_ff <= 16'd751;
        2029: data_ff <= -16'd404;
        2030: data_ff <= 16'd196;
        2031: data_ff <= -16'd77;
        2032: data_ff <= -16'd41;
        2033: data_ff <= 16'd130;
        2034: data_ff <= -16'd292;
        2035: data_ff <= 16'd562;
        2036: data_ff <= -16'd997;
        2037: data_ff <= 16'd1723;
        2038: data_ff <= -16'd3140;
        2039: data_ff <= 16'd7689;
        2040: data_ff <= 16'd30507;
        2041: data_ff <= -16'd4855;
        2042: data_ff <= 16'd2324;
        2043: data_ff <= -16'd1296;
        2044: data_ff <= 16'd733;
        2045: data_ff <= -16'd395;
        2046: data_ff <= 16'd191;
        2047: data_ff <= -16'd75;
        2048: data_ff <= -16'd40;
        2049: data_ff <= 16'd126;
        2050: data_ff <= -16'd284;
        2051: data_ff <= 16'd546;
        2052: data_ff <= -16'd969;
        2053: data_ff <= 16'd1673;
        2054: data_ff <= -16'd3046;
        2055: data_ff <= 16'd7426;
        2056: data_ff <= 16'd30638;
        2057: data_ff <= -16'd4750;
        2058: data_ff <= 16'd2269;
        2059: data_ff <= -16'd1265;
        2060: data_ff <= 16'd715;
        2061: data_ff <= -16'd385;
        2062: data_ff <= 16'd186;
        2063: data_ff <= -16'd74;
        2064: data_ff <= -16'd39;
        2065: data_ff <= 16'd122;
        2066: data_ff <= -16'd275;
        2067: data_ff <= 16'd530;
        2068: data_ff <= -16'd940;
        2069: data_ff <= 16'd1623;
        2070: data_ff <= -16'd2951;
        2071: data_ff <= 16'd7164;
        2072: data_ff <= 16'd30766;
        2073: data_ff <= -16'd4643;
        2074: data_ff <= 16'd2213;
        2075: data_ff <= -16'd1232;
        2076: data_ff <= 16'd696;
        2077: data_ff <= -16'd375;
        2078: data_ff <= 16'd182;
        2079: data_ff <= -16'd72;
        2080: data_ff <= -16'd37;
        2081: data_ff <= 16'd118;
        2082: data_ff <= -16'd267;
        2083: data_ff <= 16'd514;
        2084: data_ff <= -16'd911;
        2085: data_ff <= 16'd1572;
        2086: data_ff <= -16'd2856;
        2087: data_ff <= 16'd6904;
        2088: data_ff <= 16'd30889;
        2089: data_ff <= -16'd4532;
        2090: data_ff <= 16'd2155;
        2091: data_ff <= -16'd1199;
        2092: data_ff <= 16'd677;
        2093: data_ff <= -16'd365;
        2094: data_ff <= 16'd177;
        2095: data_ff <= -16'd70;
        2096: data_ff <= -16'd36;
        2097: data_ff <= 16'd114;
        2098: data_ff <= -16'd258;
        2099: data_ff <= 16'd497;
        2100: data_ff <= -16'd882;
        2101: data_ff <= 16'd1522;
        2102: data_ff <= -16'd2760;
        2103: data_ff <= 16'd6645;
        2104: data_ff <= 16'd31009;
        2105: data_ff <= -16'd4419;
        2106: data_ff <= 16'd2096;
        2107: data_ff <= -16'd1165;
        2108: data_ff <= 16'd658;
        2109: data_ff <= -16'd354;
        2110: data_ff <= 16'd172;
        2111: data_ff <= -16'd68;
        2112: data_ff <= -16'd35;
        2113: data_ff <= 16'd110;
        2114: data_ff <= -16'd249;
        2115: data_ff <= 16'd481;
        2116: data_ff <= -16'd853;
        2117: data_ff <= 16'd1471;
        2118: data_ff <= -16'd2664;
        2119: data_ff <= 16'd6388;
        2120: data_ff <= 16'd31125;
        2121: data_ff <= -16'd4302;
        2122: data_ff <= 16'd2035;
        2123: data_ff <= -16'd1130;
        2124: data_ff <= 16'd638;
        2125: data_ff <= -16'd343;
        2126: data_ff <= 16'd166;
        2127: data_ff <= -16'd66;
        2128: data_ff <= -16'd33;
        2129: data_ff <= 16'd107;
        2130: data_ff <= -16'd241;
        2131: data_ff <= 16'd464;
        2132: data_ff <= -16'd824;
        2133: data_ff <= 16'd1419;
        2134: data_ff <= -16'd2568;
        2135: data_ff <= 16'd6132;
        2136: data_ff <= 16'd31237;
        2137: data_ff <= -16'd4183;
        2138: data_ff <= 16'd1973;
        2139: data_ff <= -16'd1095;
        2140: data_ff <= 16'd618;
        2141: data_ff <= -16'd332;
        2142: data_ff <= 16'd161;
        2143: data_ff <= -16'd64;
        2144: data_ff <= -16'd32;
        2145: data_ff <= 16'd103;
        2146: data_ff <= -16'd232;
        2147: data_ff <= 16'd448;
        2148: data_ff <= -16'd794;
        2149: data_ff <= 16'd1368;
        2150: data_ff <= -16'd2472;
        2151: data_ff <= 16'd5878;
        2152: data_ff <= 16'd31345;
        2153: data_ff <= -16'd4060;
        2154: data_ff <= 16'd1910;
        2155: data_ff <= -16'd1059;
        2156: data_ff <= 16'd597;
        2157: data_ff <= -16'd321;
        2158: data_ff <= 16'd156;
        2159: data_ff <= -16'd62;
        2160: data_ff <= -16'd31;
        2161: data_ff <= 16'd99;
        2162: data_ff <= -16'd224;
        2163: data_ff <= 16'd431;
        2164: data_ff <= -16'd765;
        2165: data_ff <= 16'd1316;
        2166: data_ff <= -16'd2376;
        2167: data_ff <= 16'd5625;
        2168: data_ff <= 16'd31450;
        2169: data_ff <= -16'd3934;
        2170: data_ff <= 16'd1846;
        2171: data_ff <= -16'd1022;
        2172: data_ff <= 16'd576;
        2173: data_ff <= -16'd310;
        2174: data_ff <= 16'd150;
        2175: data_ff <= -16'd60;
        2176: data_ff <= -16'd29;
        2177: data_ff <= 16'd95;
        2178: data_ff <= -16'd215;
        2179: data_ff <= 16'd415;
        2180: data_ff <= -16'd735;
        2181: data_ff <= 16'd1264;
        2182: data_ff <= -16'd2279;
        2183: data_ff <= 16'd5375;
        2184: data_ff <= 16'd31550;
        2185: data_ff <= -16'd3805;
        2186: data_ff <= 16'd1781;
        2187: data_ff <= -16'd985;
        2188: data_ff <= 16'd555;
        2189: data_ff <= -16'd298;
        2190: data_ff <= 16'd145;
        2191: data_ff <= -16'd58;
        2192: data_ff <= -16'd28;
        2193: data_ff <= 16'd91;
        2194: data_ff <= -16'd206;
        2195: data_ff <= 16'd398;
        2196: data_ff <= -16'd705;
        2197: data_ff <= 16'd1213;
        2198: data_ff <= -16'd2183;
        2199: data_ff <= 16'd5125;
        2200: data_ff <= 16'd31646;
        2201: data_ff <= -16'd3673;
        2202: data_ff <= 16'd1714;
        2203: data_ff <= -16'd947;
        2204: data_ff <= 16'd533;
        2205: data_ff <= -16'd286;
        2206: data_ff <= 16'd139;
        2207: data_ff <= -16'd55;
        2208: data_ff <= -16'd27;
        2209: data_ff <= 16'd87;
        2210: data_ff <= -16'd198;
        2211: data_ff <= 16'd381;
        2212: data_ff <= -16'd676;
        2213: data_ff <= 16'd1161;
        2214: data_ff <= -16'd2086;
        2215: data_ff <= 16'd4878;
        2216: data_ff <= 16'd31738;
        2217: data_ff <= -16'd3538;
        2218: data_ff <= 16'd1646;
        2219: data_ff <= -16'd908;
        2220: data_ff <= 16'd511;
        2221: data_ff <= -16'd274;
        2222: data_ff <= 16'd133;
        2223: data_ff <= -16'd53;
        2224: data_ff <= -16'd25;
        2225: data_ff <= 16'd83;
        2226: data_ff <= -16'd189;
        2227: data_ff <= 16'd365;
        2228: data_ff <= -16'd646;
        2229: data_ff <= 16'd1108;
        2230: data_ff <= -16'd1990;
        2231: data_ff <= 16'd4633;
        2232: data_ff <= 16'd31827;
        2233: data_ff <= -16'd3400;
        2234: data_ff <= 16'd1577;
        2235: data_ff <= -16'd869;
        2236: data_ff <= 16'd488;
        2237: data_ff <= -16'd262;
        2238: data_ff <= 16'd127;
        2239: data_ff <= -16'd51;
        2240: data_ff <= -16'd24;
        2241: data_ff <= 16'd79;
        2242: data_ff <= -16'd180;
        2243: data_ff <= 16'd348;
        2244: data_ff <= -16'd616;
        2245: data_ff <= 16'd1056;
        2246: data_ff <= -16'd1893;
        2247: data_ff <= 16'd4389;
        2248: data_ff <= 16'd31911;
        2249: data_ff <= -16'd3259;
        2250: data_ff <= 16'd1507;
        2251: data_ff <= -16'd829;
        2252: data_ff <= 16'd465;
        2253: data_ff <= -16'd250;
        2254: data_ff <= 16'd121;
        2255: data_ff <= -16'd48;
        2256: data_ff <= -16'd23;
        2257: data_ff <= 16'd75;
        2258: data_ff <= -16'd172;
        2259: data_ff <= 16'd331;
        2260: data_ff <= -16'd586;
        2261: data_ff <= 16'd1004;
        2262: data_ff <= -16'd1797;
        2263: data_ff <= 16'd4147;
        2264: data_ff <= 16'd31991;
        2265: data_ff <= -16'd3115;
        2266: data_ff <= 16'd1436;
        2267: data_ff <= -16'd788;
        2268: data_ff <= 16'd442;
        2269: data_ff <= -16'd237;
        2270: data_ff <= 16'd115;
        2271: data_ff <= -16'd46;
        2272: data_ff <= -16'd22;
        2273: data_ff <= 16'd72;
        2274: data_ff <= -16'd163;
        2275: data_ff <= 16'd314;
        2276: data_ff <= -16'd556;
        2277: data_ff <= 16'd952;
        2278: data_ff <= -16'd1700;
        2279: data_ff <= 16'd3908;
        2280: data_ff <= 16'd32067;
        2281: data_ff <= -16'd2968;
        2282: data_ff <= 16'd1363;
        2283: data_ff <= -16'd747;
        2284: data_ff <= 16'd418;
        2285: data_ff <= -16'd224;
        2286: data_ff <= 16'd108;
        2287: data_ff <= -16'd43;
        2288: data_ff <= -16'd20;
        2289: data_ff <= 16'd68;
        2290: data_ff <= -16'd154;
        2291: data_ff <= 16'd298;
        2292: data_ff <= -16'd526;
        2293: data_ff <= 16'd899;
        2294: data_ff <= -16'd1604;
        2295: data_ff <= 16'd3670;
        2296: data_ff <= 16'd32138;
        2297: data_ff <= -16'd2818;
        2298: data_ff <= 16'd1290;
        2299: data_ff <= -16'd706;
        2300: data_ff <= 16'd395;
        2301: data_ff <= -16'd211;
        2302: data_ff <= 16'd102;
        2303: data_ff <= -16'd41;
        2304: data_ff <= -16'd19;
        2305: data_ff <= 16'd64;
        2306: data_ff <= -16'd146;
        2307: data_ff <= 16'd281;
        2308: data_ff <= -16'd496;
        2309: data_ff <= 16'd847;
        2310: data_ff <= -16'd1508;
        2311: data_ff <= 16'd3434;
        2312: data_ff <= 16'd32206;
        2313: data_ff <= -16'd2665;
        2314: data_ff <= 16'd1215;
        2315: data_ff <= -16'd663;
        2316: data_ff <= 16'd370;
        2317: data_ff <= -16'd198;
        2318: data_ff <= 16'd95;
        2319: data_ff <= -16'd38;
        2320: data_ff <= -16'd18;
        2321: data_ff <= 16'd60;
        2322: data_ff <= -16'd137;
        2323: data_ff <= 16'd264;
        2324: data_ff <= -16'd466;
        2325: data_ff <= 16'd795;
        2326: data_ff <= -16'd1412;
        2327: data_ff <= 16'd3201;
        2328: data_ff <= 16'd32270;
        2329: data_ff <= -16'd2509;
        2330: data_ff <= 16'd1139;
        2331: data_ff <= -16'd620;
        2332: data_ff <= 16'd346;
        2333: data_ff <= -16'd184;
        2334: data_ff <= 16'd89;
        2335: data_ff <= -16'd35;
        2336: data_ff <= -16'd17;
        2337: data_ff <= 16'd56;
        2338: data_ff <= -16'd129;
        2339: data_ff <= 16'd248;
        2340: data_ff <= -16'd436;
        2341: data_ff <= 16'd743;
        2342: data_ff <= -16'd1316;
        2343: data_ff <= 16'd2969;
        2344: data_ff <= 16'd32329;
        2345: data_ff <= -16'd2350;
        2346: data_ff <= 16'd1062;
        2347: data_ff <= -16'd577;
        2348: data_ff <= 16'd321;
        2349: data_ff <= -16'd171;
        2350: data_ff <= 16'd82;
        2351: data_ff <= -16'd33;
        2352: data_ff <= -16'd16;
        2353: data_ff <= 16'd53;
        2354: data_ff <= -16'd120;
        2355: data_ff <= 16'd231;
        2356: data_ff <= -16'd406;
        2357: data_ff <= 16'd691;
        2358: data_ff <= -16'd1221;
        2359: data_ff <= 16'd2740;
        2360: data_ff <= 16'd32384;
        2361: data_ff <= -16'd2189;
        2362: data_ff <= 16'd985;
        2363: data_ff <= -16'd533;
        2364: data_ff <= 16'd296;
        2365: data_ff <= -16'd157;
        2366: data_ff <= 16'd75;
        2367: data_ff <= -16'd30;
        2368: data_ff <= -16'd14;
        2369: data_ff <= 16'd49;
        2370: data_ff <= -16'd111;
        2371: data_ff <= 16'd214;
        2372: data_ff <= -16'd377;
        2373: data_ff <= 16'd639;
        2374: data_ff <= -16'd1126;
        2375: data_ff <= 16'd2513;
        2376: data_ff <= 16'd32435;
        2377: data_ff <= -16'd2024;
        2378: data_ff <= 16'd906;
        2379: data_ff <= -16'd489;
        2380: data_ff <= 16'd270;
        2381: data_ff <= -16'd143;
        2382: data_ff <= 16'd68;
        2383: data_ff <= -16'd27;
        2384: data_ff <= -16'd13;
        2385: data_ff <= 16'd45;
        2386: data_ff <= -16'd103;
        2387: data_ff <= 16'd198;
        2388: data_ff <= -16'd347;
        2389: data_ff <= 16'd587;
        2390: data_ff <= -16'd1031;
        2391: data_ff <= 16'd2288;
        2392: data_ff <= 16'd32482;
        2393: data_ff <= -16'd1856;
        2394: data_ff <= 16'd826;
        2395: data_ff <= -16'd444;
        2396: data_ff <= 16'd244;
        2397: data_ff <= -16'd129;
        2398: data_ff <= 16'd61;
        2399: data_ff <= -16'd24;
        2400: data_ff <= -16'd12;
        2401: data_ff <= 16'd41;
        2402: data_ff <= -16'd95;
        2403: data_ff <= 16'd181;
        2404: data_ff <= -16'd317;
        2405: data_ff <= 16'd535;
        2406: data_ff <= -16'd936;
        2407: data_ff <= 16'd2065;
        2408: data_ff <= 16'd32525;
        2409: data_ff <= -16'd1686;
        2410: data_ff <= 16'd745;
        2411: data_ff <= -16'd399;
        2412: data_ff <= 16'd218;
        2413: data_ff <= -16'd114;
        2414: data_ff <= 16'd54;
        2415: data_ff <= -16'd21;
        2416: data_ff <= -16'd11;
        2417: data_ff <= 16'd38;
        2418: data_ff <= -16'd86;
        2419: data_ff <= 16'd165;
        2420: data_ff <= -16'd287;
        2421: data_ff <= 16'd483;
        2422: data_ff <= -16'd842;
        2423: data_ff <= 16'd1845;
        2424: data_ff <= 16'd32563;
        2425: data_ff <= -16'd1513;
        2426: data_ff <= 16'd664;
        2427: data_ff <= -16'd353;
        2428: data_ff <= 16'd192;
        2429: data_ff <= -16'd100;
        2430: data_ff <= 16'd47;
        2431: data_ff <= -16'd18;
        2432: data_ff <= -16'd10;
        2433: data_ff <= 16'd34;
        2434: data_ff <= -16'd78;
        2435: data_ff <= 16'd148;
        2436: data_ff <= -16'd258;
        2437: data_ff <= 16'd432;
        2438: data_ff <= -16'd749;
        2439: data_ff <= 16'd1627;
        2440: data_ff <= 16'd32597;
        2441: data_ff <= -16'd1337;
        2442: data_ff <= 16'd581;
        2443: data_ff <= -16'd306;
        2444: data_ff <= 16'd165;
        2445: data_ff <= -16'd85;
        2446: data_ff <= 16'd40;
        2447: data_ff <= -16'd15;
        2448: data_ff <= -16'd9;
        2449: data_ff <= 16'd31;
        2450: data_ff <= -16'd69;
        2451: data_ff <= 16'd132;
        2452: data_ff <= -16'd228;
        2453: data_ff <= 16'd381;
        2454: data_ff <= -16'd656;
        2455: data_ff <= 16'd1412;
        2456: data_ff <= 16'd32627;
        2457: data_ff <= -16'd1158;
        2458: data_ff <= 16'd498;
        2459: data_ff <= -16'd260;
        2460: data_ff <= 16'd139;
        2461: data_ff <= -16'd71;
        2462: data_ff <= 16'd32;
        2463: data_ff <= -16'd12;
        2464: data_ff <= -16'd8;
        2465: data_ff <= 16'd27;
        2466: data_ff <= -16'd61;
        2467: data_ff <= 16'd116;
        2468: data_ff <= -16'd199;
        2469: data_ff <= 16'd330;
        2470: data_ff <= -16'd563;
        2471: data_ff <= 16'd1199;
        2472: data_ff <= 16'd32653;
        2473: data_ff <= -16'd976;
        2474: data_ff <= 16'd413;
        2475: data_ff <= -16'd212;
        2476: data_ff <= 16'd111;
        2477: data_ff <= -16'd56;
        2478: data_ff <= 16'd25;
        2479: data_ff <= -16'd9;
        2480: data_ff <= -16'd7;
        2481: data_ff <= 16'd23;
        2482: data_ff <= -16'd53;
        2483: data_ff <= 16'd100;
        2484: data_ff <= -16'd170;
        2485: data_ff <= 16'd279;
        2486: data_ff <= -16'd471;
        2487: data_ff <= 16'd988;
        2488: data_ff <= 16'd32674;
        2489: data_ff <= -16'd791;
        2490: data_ff <= 16'd328;
        2491: data_ff <= -16'd165;
        2492: data_ff <= 16'd84;
        2493: data_ff <= -16'd41;
        2494: data_ff <= 16'd17;
        2495: data_ff <= -16'd6;
        2496: data_ff <= -16'd6;
        2497: data_ff <= 16'd20;
        2498: data_ff <= -16'd45;
        2499: data_ff <= 16'd83;
        2500: data_ff <= -16'd141;
        2501: data_ff <= 16'd228;
        2502: data_ff <= -16'd380;
        2503: data_ff <= 16'd780;
        2504: data_ff <= 16'd32691;
        2505: data_ff <= -16'd604;
        2506: data_ff <= 16'd242;
        2507: data_ff <= -16'd117;
        2508: data_ff <= 16'd57;
        2509: data_ff <= -16'd25;
        2510: data_ff <= 16'd10;
        2511: data_ff <= -16'd3;
        2512: data_ff <= -16'd5;
        2513: data_ff <= 16'd16;
        2514: data_ff <= -16'd37;
        2515: data_ff <= 16'd67;
        2516: data_ff <= -16'd112;
        2517: data_ff <= 16'd178;
        2518: data_ff <= -16'd289;
        2519: data_ff <= 16'd574;
        2520: data_ff <= 16'd32704;
        2521: data_ff <= -16'd414;
        2522: data_ff <= 16'd155;
        2523: data_ff <= -16'd68;
        2524: data_ff <= 16'd29;
        2525: data_ff <= -16'd10;
        2526: data_ff <= 16'd2;
        2527: data_ff <= 16'd0;
        2528: data_ff <= -16'd4;
        2529: data_ff <= 16'd13;
        2530: data_ff <= -16'd29;
        2531: data_ff <= 16'd52;
        2532: data_ff <= -16'd83;
        2533: data_ff <= 16'd128;
        2534: data_ff <= -16'd198;
        2535: data_ff <= 16'd371;
        2536: data_ff <= 16'd32712;
        2537: data_ff <= -16'd222;
        2538: data_ff <= 16'd68;
        2539: data_ff <= -16'd20;
        2540: data_ff <= 16'd1;
        2541: data_ff <= 16'd4;
        2542: data_ff <= -16'd5;
        2543: data_ff <= 16'd3;
        2544: data_ff <= -16'd3;
        2545: data_ff <= 16'd10;
        2546: data_ff <= -16'd21;
        2547: data_ff <= 16'd36;
        2548: data_ff <= -16'd55;
        2549: data_ff <= 16'd78;
        2550: data_ff <= -16'd109;
        2551: data_ff <= 16'd171;
        2552: data_ff <= 16'd32717;
        2553: data_ff <= -16'd26;
        2554: data_ff <= -16'd20;
        2555: data_ff <= 16'd29;
        2556: data_ff <= -16'd26;
        2557: data_ff <= 16'd20;
        2558: data_ff <= -16'd13;
        2559: data_ff <= 16'd6;
        default: data_ff <= 0;
    endcase
end
endmodule
