
module rom_firbank_441_480(
    input clk,
    input [10:0] addr,
    output [23:0] data);
reg [23:0] data_ff;
assign data = data_ff;
always @(posedge clk) begin
    case(addr)
        0: data_ff <= 24'd43559;
        1: data_ff <= -24'd27408;
        2: data_ff <= 24'd19328;
        3: data_ff <= -24'd13322;
        4: data_ff <= 24'd8607;
        5: data_ff <= -24'd5089;
        6: data_ff <= 24'd2693;
        7: data_ff <= -24'd1241;
        8: data_ff <= 24'd476;
        9: data_ff <= -24'd141;
        10: data_ff <= 24'd25;
        11: data_ff <= -24'd1;
        12: data_ff <= 24'd94619;
        13: data_ff <= -24'd49936;
        14: data_ff <= 24'd31583;
        15: data_ff <= -24'd20206;
        16: data_ff <= 24'd12364;
        17: data_ff <= -24'd7015;
        18: data_ff <= 24'd3595;
        19: data_ff <= -24'd1613;
        20: data_ff <= 24'd607;
        21: data_ff <= -24'd176;
        22: data_ff <= 24'd31;
        23: data_ff <= -24'd1;
        24: data_ff <= 24'd146342;
        25: data_ff <= -24'd72632;
        26: data_ff <= 24'd43915;
        27: data_ff <= -24'd27132;
        28: data_ff <= 24'd16146;
        29: data_ff <= -24'd8955;
        30: data_ff <= 24'd4504;
        31: data_ff <= -24'd1990;
        32: data_ff <= 24'd739;
        33: data_ff <= -24'd212;
        34: data_ff <= 24'd37;
        35: data_ff <= -24'd1;
        36: data_ff <= 24'd198719;
        37: data_ff <= -24'd95488;
        38: data_ff <= 24'd56319;
        39: data_ff <= -24'd34098;
        40: data_ff <= 24'd19952;
        41: data_ff <= -24'd10909;
        42: data_ff <= 24'd5420;
        43: data_ff <= -24'd2371;
        44: data_ff <= 24'd872;
        45: data_ff <= -24'd249;
        46: data_ff <= 24'd44;
        47: data_ff <= -24'd2;
        48: data_ff <= 24'd251742;
        49: data_ff <= -24'd118497;
        50: data_ff <= 24'd68790;
        51: data_ff <= -24'd41102;
        52: data_ff <= 24'd23780;
        53: data_ff <= -24'd12876;
        54: data_ff <= 24'd6344;
        55: data_ff <= -24'd2755;
        56: data_ff <= 24'd1008;
        57: data_ff <= -24'd286;
        58: data_ff <= 24'd50;
        59: data_ff <= -24'd2;
        60: data_ff <= 24'd305404;
        61: data_ff <= -24'd141651;
        62: data_ff <= 24'd81325;
        63: data_ff <= -24'd48141;
        64: data_ff <= 24'd27629;
        65: data_ff <= -24'd14855;
        66: data_ff <= 24'd7274;
        67: data_ff <= -24'd3142;
        68: data_ff <= 24'd1144;
        69: data_ff <= -24'd324;
        70: data_ff <= 24'd57;
        71: data_ff <= -24'd2;
        72: data_ff <= 24'd359697;
        73: data_ff <= -24'd164943;
        74: data_ff <= 24'd93919;
        75: data_ff <= -24'd55212;
        76: data_ff <= 24'd31498;
        77: data_ff <= -24'd16846;
        78: data_ff <= 24'd8211;
        79: data_ff <= -24'd3533;
        80: data_ff <= 24'd1283;
        81: data_ff <= -24'd363;
        82: data_ff <= 24'd64;
        83: data_ff <= -24'd2;
        84: data_ff <= 24'd414612;
        85: data_ff <= -24'd188365;
        86: data_ff <= 24'd106568;
        87: data_ff <= -24'd62313;
        88: data_ff <= 24'd35384;
        89: data_ff <= -24'd18848;
        90: data_ff <= 24'd9154;
        91: data_ff <= -24'd3927;
        92: data_ff <= 24'd1422;
        93: data_ff <= -24'd402;
        94: data_ff <= 24'd71;
        95: data_ff <= -24'd3;
        96: data_ff <= 24'd470140;
        97: data_ff <= -24'd211910;
        98: data_ff <= 24'd119266;
        99: data_ff <= -24'd69441;
        100: data_ff <= 24'd39287;
        101: data_ff <= -24'd20860;
        102: data_ff <= 24'd10103;
        103: data_ff <= -24'd4324;
        104: data_ff <= 24'd1563;
        105: data_ff <= -24'd441;
        106: data_ff <= 24'd78;
        107: data_ff <= -24'd3;
        108: data_ff <= 24'd526274;
        109: data_ff <= -24'd235568;
        110: data_ff <= 24'd132009;
        111: data_ff <= -24'd76594;
        112: data_ff <= 24'd43204;
        113: data_ff <= -24'd22881;
        114: data_ff <= 24'd11058;
        115: data_ff <= -24'd4724;
        116: data_ff <= 24'd1706;
        117: data_ff <= -24'd481;
        118: data_ff <= 24'd85;
        119: data_ff <= -24'd3;
        120: data_ff <= 24'd583002;
        121: data_ff <= -24'd259333;
        122: data_ff <= 24'd144792;
        123: data_ff <= -24'd83768;
        124: data_ff <= 24'd47136;
        125: data_ff <= -24'd24910;
        126: data_ff <= 24'd12017;
        127: data_ff <= -24'd5127;
        128: data_ff <= 24'd1850;
        129: data_ff <= -24'd522;
        130: data_ff <= 24'd93;
        131: data_ff <= -24'd4;
        132: data_ff <= 24'd640318;
        133: data_ff <= -24'd283195;
        134: data_ff <= 24'd157611;
        135: data_ff <= -24'd90961;
        136: data_ff <= 24'd51079;
        137: data_ff <= -24'd26948;
        138: data_ff <= 24'd12982;
        139: data_ff <= -24'd5532;
        140: data_ff <= 24'd1995;
        141: data_ff <= -24'd563;
        142: data_ff <= 24'd100;
        143: data_ff <= -24'd4;
        144: data_ff <= 24'd698211;
        145: data_ff <= -24'd307147;
        146: data_ff <= 24'd170461;
        147: data_ff <= -24'd98171;
        148: data_ff <= 24'd55033;
        149: data_ff <= -24'd28993;
        150: data_ff <= 24'd13950;
        151: data_ff <= -24'd5940;
        152: data_ff <= 24'd2141;
        153: data_ff <= -24'd604;
        154: data_ff <= 24'd108;
        155: data_ff <= -24'd4;
        156: data_ff <= 24'd756671;
        157: data_ff <= -24'd331181;
        158: data_ff <= 24'd183337;
        159: data_ff <= -24'd105395;
        160: data_ff <= 24'd58997;
        161: data_ff <= -24'd31043;
        162: data_ff <= 24'd14923;
        163: data_ff <= -24'd6350;
        164: data_ff <= 24'd2288;
        165: data_ff <= -24'd646;
        166: data_ff <= 24'd116;
        167: data_ff <= -24'd5;
        168: data_ff <= 24'd815689;
        169: data_ff <= -24'd355287;
        170: data_ff <= 24'd196234;
        171: data_ff <= -24'd112629;
        172: data_ff <= 24'd62967;
        173: data_ff <= -24'd33100;
        174: data_ff <= 24'd15900;
        175: data_ff <= -24'd6762;
        176: data_ff <= 24'd2436;
        177: data_ff <= -24'd689;
        178: data_ff <= 24'd124;
        179: data_ff <= -24'd5;
        180: data_ff <= 24'd875255;
        181: data_ff <= -24'd379458;
        182: data_ff <= 24'd209147;
        183: data_ff <= -24'd119871;
        184: data_ff <= 24'd66944;
        185: data_ff <= -24'd35161;
        186: data_ff <= 24'd16880;
        187: data_ff <= -24'd7177;
        188: data_ff <= 24'd2586;
        189: data_ff <= -24'd731;
        190: data_ff <= 24'd132;
        191: data_ff <= -24'd5;
        192: data_ff <= 24'd935359;
        193: data_ff <= -24'd403684;
        194: data_ff <= 24'd222071;
        195: data_ff <= -24'd127118;
        196: data_ff <= 24'd70925;
        197: data_ff <= -24'd37226;
        198: data_ff <= 24'd17862;
        199: data_ff <= -24'd7593;
        200: data_ff <= 24'd2736;
        201: data_ff <= -24'd775;
        202: data_ff <= 24'd140;
        203: data_ff <= -24'd6;
        204: data_ff <= 24'd995990;
        205: data_ff <= -24'd427958;
        206: data_ff <= 24'd235002;
        207: data_ff <= -24'd134367;
        208: data_ff <= 24'd74908;
        209: data_ff <= -24'd39293;
        210: data_ff <= 24'd18848;
        211: data_ff <= -24'd8011;
        212: data_ff <= 24'd2888;
        213: data_ff <= -24'd818;
        214: data_ff <= 24'd149;
        215: data_ff <= -24'd6;
        216: data_ff <= 24'd1057138;
        217: data_ff <= -24'd452269;
        218: data_ff <= 24'd247933;
        219: data_ff <= -24'd141616;
        220: data_ff <= 24'd78893;
        221: data_ff <= -24'd41364;
        222: data_ff <= 24'd19835;
        223: data_ff <= -24'd8430;
        224: data_ff <= 24'd3040;
        225: data_ff <= -24'd862;
        226: data_ff <= 24'd157;
        227: data_ff <= -24'd7;
        228: data_ff <= 24'd1118792;
        229: data_ff <= -24'd476609;
        230: data_ff <= 24'd260861;
        231: data_ff <= -24'd148861;
        232: data_ff <= 24'd82878;
        233: data_ff <= -24'd43435;
        234: data_ff <= 24'd20824;
        235: data_ff <= -24'd8851;
        236: data_ff <= 24'd3193;
        237: data_ff <= -24'd907;
        238: data_ff <= 24'd166;
        239: data_ff <= -24'd7;
        240: data_ff <= 24'd1180942;
        241: data_ff <= -24'd500970;
        242: data_ff <= 24'd273779;
        243: data_ff <= -24'd156099;
        244: data_ff <= 24'd86860;
        245: data_ff <= -24'd45507;
        246: data_ff <= 24'd21815;
        247: data_ff <= -24'd9273;
        248: data_ff <= 24'd3347;
        249: data_ff <= -24'd952;
        250: data_ff <= 24'd175;
        251: data_ff <= -24'd7;
        252: data_ff <= 24'd1243575;
        253: data_ff <= -24'd525342;
        254: data_ff <= 24'd286683;
        255: data_ff <= -24'd163328;
        256: data_ff <= 24'd90839;
        257: data_ff <= -24'd47579;
        258: data_ff <= 24'd22806;
        259: data_ff <= -24'd9696;
        260: data_ff <= 24'd3502;
        261: data_ff <= -24'd997;
        262: data_ff <= 24'd184;
        263: data_ff <= -24'd8;
        264: data_ff <= 24'd1306682;
        265: data_ff <= -24'd549715;
        266: data_ff <= 24'd299568;
        267: data_ff <= -24'd170545;
        268: data_ff <= 24'd94813;
        269: data_ff <= -24'd49649;
        270: data_ff <= 24'd23798;
        271: data_ff <= -24'd10120;
        272: data_ff <= 24'd3657;
        273: data_ff <= -24'd1042;
        274: data_ff <= 24'd193;
        275: data_ff <= -24'd8;
        276: data_ff <= 24'd1370250;
        277: data_ff <= -24'd574082;
        278: data_ff <= 24'd312428;
        279: data_ff <= -24'd177746;
        280: data_ff <= 24'd98779;
        281: data_ff <= -24'd51717;
        282: data_ff <= 24'd24790;
        283: data_ff <= -24'd10545;
        284: data_ff <= 24'd3813;
        285: data_ff <= -24'd1088;
        286: data_ff <= 24'd202;
        287: data_ff <= -24'd9;
        288: data_ff <= 24'd1434267;
        289: data_ff <= -24'd598431;
        290: data_ff <= 24'd325258;
        291: data_ff <= -24'd184929;
        292: data_ff <= 24'd102737;
        293: data_ff <= -24'd53783;
        294: data_ff <= 24'd25782;
        295: data_ff <= -24'd10970;
        296: data_ff <= 24'd3969;
        297: data_ff <= -24'd1134;
        298: data_ff <= 24'd212;
        299: data_ff <= -24'd9;
        300: data_ff <= 24'd1498724;
        301: data_ff <= -24'd622755;
        302: data_ff <= 24'd338053;
        303: data_ff <= -24'd192090;
        304: data_ff <= 24'd106684;
        305: data_ff <= -24'd55844;
        306: data_ff <= 24'd26773;
        307: data_ff <= -24'd11396;
        308: data_ff <= 24'd4126;
        309: data_ff <= -24'd1181;
        310: data_ff <= 24'd221;
        311: data_ff <= -24'd10;
        312: data_ff <= 24'd1563606;
        313: data_ff <= -24'd647043;
        314: data_ff <= 24'd350808;
        315: data_ff <= -24'd199227;
        316: data_ff <= 24'd110620;
        317: data_ff <= -24'd57901;
        318: data_ff <= 24'd27763;
        319: data_ff <= -24'd11822;
        320: data_ff <= 24'd4283;
        321: data_ff <= -24'd1227;
        322: data_ff <= 24'd231;
        323: data_ff <= -24'd10;
        324: data_ff <= 24'd1628903;
        325: data_ff <= -24'd671287;
        326: data_ff <= 24'd363516;
        327: data_ff <= -24'd206336;
        328: data_ff <= 24'd114541;
        329: data_ff <= -24'd59952;
        330: data_ff <= 24'd28751;
        331: data_ff <= -24'd12247;
        332: data_ff <= 24'd4440;
        333: data_ff <= -24'd1274;
        334: data_ff <= 24'd240;
        335: data_ff <= -24'd11;
        336: data_ff <= 24'd1694601;
        337: data_ff <= -24'd695476;
        338: data_ff <= 24'd376174;
        339: data_ff <= -24'd213415;
        340: data_ff <= 24'd118447;
        341: data_ff <= -24'd61997;
        342: data_ff <= 24'd29738;
        343: data_ff <= -24'd12673;
        344: data_ff <= 24'd4598;
        345: data_ff <= -24'd1321;
        346: data_ff <= 24'd250;
        347: data_ff <= -24'd12;
        348: data_ff <= 24'd1760690;
        349: data_ff <= -24'd719600;
        350: data_ff <= 24'd388775;
        351: data_ff <= -24'd220460;
        352: data_ff <= 24'd122336;
        353: data_ff <= -24'd64035;
        354: data_ff <= 24'd30722;
        355: data_ff <= -24'd13098;
        356: data_ff <= 24'd4756;
        357: data_ff <= -24'd1369;
        358: data_ff <= 24'd260;
        359: data_ff <= -24'd12;
        360: data_ff <= 24'd1827155;
        361: data_ff <= -24'd743651;
        362: data_ff <= 24'd401314;
        363: data_ff <= -24'd227468;
        364: data_ff <= 24'd126207;
        365: data_ff <= -24'd66064;
        366: data_ff <= 24'd31702;
        367: data_ff <= -24'd13522;
        368: data_ff <= 24'd4914;
        369: data_ff <= -24'd1416;
        370: data_ff <= 24'd270;
        371: data_ff <= -24'd13;
        372: data_ff <= 24'd1893985;
        373: data_ff <= -24'd767618;
        374: data_ff <= 24'd413785;
        375: data_ff <= -24'd234436;
        376: data_ff <= 24'd130056;
        377: data_ff <= -24'd68083;
        378: data_ff <= 24'd32680;
        379: data_ff <= -24'd13946;
        380: data_ff <= 24'd5072;
        381: data_ff <= -24'd1464;
        382: data_ff <= 24'd280;
        383: data_ff <= -24'd14;
        384: data_ff <= 24'd1961166;
        385: data_ff <= -24'd791492;
        386: data_ff <= 24'd426184;
        387: data_ff <= -24'd241362;
        388: data_ff <= 24'd133883;
        389: data_ff <= -24'd70093;
        390: data_ff <= 24'd33654;
        391: data_ff <= -24'd14368;
        392: data_ff <= 24'd5230;
        393: data_ff <= -24'd1512;
        394: data_ff <= 24'd290;
        395: data_ff <= -24'd14;
        396: data_ff <= 24'd2028686;
        397: data_ff <= -24'd815263;
        398: data_ff <= 24'd438506;
        399: data_ff <= -24'd248242;
        400: data_ff <= 24'd137687;
        401: data_ff <= -24'd72092;
        402: data_ff <= 24'd34623;
        403: data_ff <= -24'd14790;
        404: data_ff <= 24'd5388;
        405: data_ff <= -24'd1560;
        406: data_ff <= 24'd300;
        407: data_ff <= -24'd15;
        408: data_ff <= 24'd2096532;
        409: data_ff <= -24'd838920;
        410: data_ff <= 24'd450743;
        411: data_ff <= -24'd255072;
        412: data_ff <= 24'd141464;
        413: data_ff <= -24'd74078;
        414: data_ff <= 24'd35588;
        415: data_ff <= -24'd15210;
        416: data_ff <= 24'd5546;
        417: data_ff <= -24'd1608;
        418: data_ff <= 24'd311;
        419: data_ff <= -24'd16;
        420: data_ff <= 24'd2164689;
        421: data_ff <= -24'd862455;
        422: data_ff <= 24'd462892;
        423: data_ff <= -24'd261851;
        424: data_ff <= 24'd145214;
        425: data_ff <= -24'd76052;
        426: data_ff <= 24'd36548;
        427: data_ff <= -24'd15629;
        428: data_ff <= 24'd5703;
        429: data_ff <= -24'd1656;
        430: data_ff <= 24'd321;
        431: data_ff <= -24'd17;
        432: data_ff <= 24'd2233146;
        433: data_ff <= -24'd885856;
        434: data_ff <= 24'd474946;
        435: data_ff <= -24'd268574;
        436: data_ff <= 24'd148935;
        437: data_ff <= -24'd78012;
        438: data_ff <= 24'd37502;
        439: data_ff <= -24'd16045;
        440: data_ff <= 24'd5861;
        441: data_ff <= -24'd1704;
        442: data_ff <= 24'd332;
        443: data_ff <= -24'd17;
        444: data_ff <= 24'd2301888;
        445: data_ff <= -24'd909115;
        446: data_ff <= 24'd486900;
        447: data_ff <= -24'd275239;
        448: data_ff <= 24'd152625;
        449: data_ff <= -24'd79957;
        450: data_ff <= 24'd38450;
        451: data_ff <= -24'd16460;
        452: data_ff <= 24'd6018;
        453: data_ff <= -24'd1752;
        454: data_ff <= 24'd342;
        455: data_ff <= -24'd18;
        456: data_ff <= 24'd2370902;
        457: data_ff <= -24'd932221;
        458: data_ff <= 24'd498749;
        459: data_ff <= -24'd281843;
        460: data_ff <= 24'd156282;
        461: data_ff <= -24'd81887;
        462: data_ff <= 24'd39392;
        463: data_ff <= -24'd16873;
        464: data_ff <= 24'd6174;
        465: data_ff <= -24'd1801;
        466: data_ff <= 24'd353;
        467: data_ff <= -24'd19;
        468: data_ff <= 24'd2440174;
        469: data_ff <= -24'd955163;
        470: data_ff <= 24'd510488;
        471: data_ff <= -24'd288382;
        472: data_ff <= 24'd159904;
        473: data_ff <= -24'd83800;
        474: data_ff <= 24'd40326;
        475: data_ff <= -24'd17283;
        476: data_ff <= 24'd6330;
        477: data_ff <= -24'd1849;
        478: data_ff <= 24'd364;
        479: data_ff <= -24'd20;
        480: data_ff <= 24'd2509690;
        481: data_ff <= -24'd977932;
        482: data_ff <= 24'd522110;
        483: data_ff <= -24'd294854;
        484: data_ff <= 24'd163490;
        485: data_ff <= -24'd85695;
        486: data_ff <= 24'd41253;
        487: data_ff <= -24'd17691;
        488: data_ff <= 24'd6485;
        489: data_ff <= -24'd1897;
        490: data_ff <= 24'd374;
        491: data_ff <= -24'd21;
        492: data_ff <= 24'd2579436;
        493: data_ff <= -24'd1000518;
        494: data_ff <= 24'd533611;
        495: data_ff <= -24'd301255;
        496: data_ff <= 24'd167039;
        497: data_ff <= -24'd87572;
        498: data_ff <= 24'd42173;
        499: data_ff <= -24'd18095;
        500: data_ff <= 24'd6639;
        501: data_ff <= -24'd1945;
        502: data_ff <= 24'd385;
        503: data_ff <= -24'd22;
        504: data_ff <= 24'd2649399;
        505: data_ff <= -24'd1022911;
        506: data_ff <= 24'd544985;
        507: data_ff <= -24'd307582;
        508: data_ff <= 24'd170548;
        509: data_ff <= -24'd89429;
        510: data_ff <= 24'd43083;
        511: data_ff <= -24'd18497;
        512: data_ff <= 24'd6793;
        513: data_ff <= -24'd1993;
        514: data_ff <= 24'd396;
        515: data_ff <= -24'd23;
        516: data_ff <= 24'd2719563;
        517: data_ff <= -24'd1045100;
        518: data_ff <= 24'd556227;
        519: data_ff <= -24'd313832;
        520: data_ff <= 24'd174015;
        521: data_ff <= -24'd91266;
        522: data_ff <= 24'd43985;
        523: data_ff <= -24'd18896;
        524: data_ff <= 24'd6946;
        525: data_ff <= -24'd2041;
        526: data_ff <= 24'd407;
        527: data_ff <= -24'd24;
        528: data_ff <= 24'd2789915;
        529: data_ff <= -24'd1067075;
        530: data_ff <= 24'd567331;
        531: data_ff <= -24'd320003;
        532: data_ff <= 24'd177439;
        533: data_ff <= -24'd93082;
        534: data_ff <= 24'd44878;
        535: data_ff <= -24'd19291;
        536: data_ff <= 24'd7097;
        537: data_ff <= -24'd2089;
        538: data_ff <= 24'd418;
        539: data_ff <= -24'd25;
        540: data_ff <= 24'd2860440;
        541: data_ff <= -24'd1088826;
        542: data_ff <= 24'd578292;
        543: data_ff <= -24'd326091;
        544: data_ff <= 24'd180818;
        545: data_ff <= -24'd94875;
        546: data_ff <= 24'd45761;
        547: data_ff <= -24'd19683;
        548: data_ff <= 24'd7248;
        549: data_ff <= -24'd2136;
        550: data_ff <= 24'd429;
        551: data_ff <= -24'd26;
        552: data_ff <= 24'd2931123;
        553: data_ff <= -24'd1110343;
        554: data_ff <= 24'd589105;
        555: data_ff <= -24'd332092;
        556: data_ff <= 24'd184151;
        557: data_ff <= -24'd96646;
        558: data_ff <= 24'd46634;
        559: data_ff <= -24'd20070;
        560: data_ff <= 24'd7398;
        561: data_ff <= -24'd2184;
        562: data_ff <= 24'd440;
        563: data_ff <= -24'd27;
        564: data_ff <= 24'd3001951;
        565: data_ff <= -24'd1131616;
        566: data_ff <= 24'd599763;
        567: data_ff <= -24'd338005;
        568: data_ff <= 24'd187436;
        569: data_ff <= -24'd98392;
        570: data_ff <= 24'd47496;
        571: data_ff <= -24'd20454;
        572: data_ff <= 24'd7546;
        573: data_ff <= -24'd2231;
        574: data_ff <= 24'd451;
        575: data_ff <= -24'd28;
        576: data_ff <= 24'd3072908;
        577: data_ff <= -24'd1152634;
        578: data_ff <= 24'd610263;
        579: data_ff <= -24'd343826;
        580: data_ff <= 24'd190670;
        581: data_ff <= -24'd100113;
        582: data_ff <= 24'd48346;
        583: data_ff <= -24'd20833;
        584: data_ff <= 24'd7693;
        585: data_ff <= -24'd2278;
        586: data_ff <= 24'd462;
        587: data_ff <= -24'd29;
        588: data_ff <= 24'd3143980;
        589: data_ff <= -24'd1173388;
        590: data_ff <= 24'd620598;
        591: data_ff <= -24'd349552;
        592: data_ff <= 24'd193853;
        593: data_ff <= -24'd101808;
        594: data_ff <= 24'd49185;
        595: data_ff <= -24'd21208;
        596: data_ff <= 24'd7839;
        597: data_ff <= -24'd2324;
        598: data_ff <= 24'd473;
        599: data_ff <= -24'd30;
        600: data_ff <= 24'd3215152;
        601: data_ff <= -24'd1193866;
        602: data_ff <= 24'd630764;
        603: data_ff <= -24'd355180;
        604: data_ff <= 24'd196982;
        605: data_ff <= -24'd103477;
        606: data_ff <= 24'd50012;
        607: data_ff <= -24'd21578;
        608: data_ff <= 24'd7984;
        609: data_ff <= -24'd2371;
        610: data_ff <= 24'd484;
        611: data_ff <= -24'd31;
        612: data_ff <= 24'd3286409;
        613: data_ff <= -24'd1214060;
        614: data_ff <= 24'd640754;
        615: data_ff <= -24'd360707;
        616: data_ff <= 24'd200057;
        617: data_ff <= -24'd105117;
        618: data_ff <= 24'd50827;
        619: data_ff <= -24'd21944;
        620: data_ff <= 24'd8126;
        621: data_ff <= -24'd2417;
        622: data_ff <= 24'd495;
        623: data_ff <= -24'd32;
        624: data_ff <= 24'd3357735;
        625: data_ff <= -24'd1233958;
        626: data_ff <= 24'd650565;
        627: data_ff <= -24'd366130;
        628: data_ff <= 24'd203074;
        629: data_ff <= -24'd106729;
        630: data_ff <= 24'd51628;
        631: data_ff <= -24'd22304;
        632: data_ff <= 24'd8268;
        633: data_ff <= -24'd2463;
        634: data_ff <= 24'd506;
        635: data_ff <= -24'd33;
        636: data_ff <= 24'd3429117;
        637: data_ff <= -24'd1253552;
        638: data_ff <= 24'd660190;
        639: data_ff <= -24'd371447;
        640: data_ff <= 24'd206033;
        641: data_ff <= -24'd108312;
        642: data_ff <= 24'd52416;
        643: data_ff <= -24'd22659;
        644: data_ff <= 24'd8407;
        645: data_ff <= -24'd2508;
        646: data_ff <= 24'd516;
        647: data_ff <= -24'd34;
        648: data_ff <= 24'd3500538;
        649: data_ff <= -24'd1272829;
        650: data_ff <= 24'd669625;
        651: data_ff <= -24'd376654;
        652: data_ff <= 24'd208933;
        653: data_ff <= -24'd109863;
        654: data_ff <= 24'd53190;
        655: data_ff <= -24'd23008;
        656: data_ff <= 24'd8545;
        657: data_ff <= -24'd2553;
        658: data_ff <= 24'd527;
        659: data_ff <= -24'd36;
        660: data_ff <= 24'd3571984;
        661: data_ff <= -24'd1291781;
        662: data_ff <= 24'd678864;
        663: data_ff <= -24'd381748;
        664: data_ff <= 24'd211770;
        665: data_ff <= -24'd111384;
        666: data_ff <= 24'd53949;
        667: data_ff <= -24'd23351;
        668: data_ff <= 24'd8680;
        669: data_ff <= -24'd2597;
        670: data_ff <= 24'd538;
        671: data_ff <= -24'd37;
        672: data_ff <= 24'd3643439;
        673: data_ff <= -24'd1310397;
        674: data_ff <= 24'd687902;
        675: data_ff <= -24'd386727;
        676: data_ff <= 24'd214544;
        677: data_ff <= -24'd112872;
        678: data_ff <= 24'd54694;
        679: data_ff <= -24'd23689;
        680: data_ff <= 24'd8814;
        681: data_ff <= -24'd2641;
        682: data_ff <= 24'd549;
        683: data_ff <= -24'd38;
        684: data_ff <= 24'd3714888;
        685: data_ff <= -24'd1328668;
        686: data_ff <= 24'd696735;
        687: data_ff <= -24'd391588;
        688: data_ff <= 24'd217254;
        689: data_ff <= -24'd114327;
        690: data_ff <= 24'd55423;
        691: data_ff <= -24'd24020;
        692: data_ff <= 24'd8946;
        693: data_ff <= -24'd2685;
        694: data_ff <= 24'd560;
        695: data_ff <= -24'd39;
        696: data_ff <= 24'd3786316;
        697: data_ff <= -24'd1346582;
        698: data_ff <= 24'd705358;
        699: data_ff <= -24'd396328;
        700: data_ff <= 24'd219896;
        701: data_ff <= -24'd115748;
        702: data_ff <= 24'd56136;
        703: data_ff <= -24'd24345;
        704: data_ff <= 24'd9076;
        705: data_ff <= -24'd2728;
        706: data_ff <= 24'd571;
        707: data_ff <= -24'd41;
        708: data_ff <= 24'd3857707;
        709: data_ff <= -24'd1364131;
        710: data_ff <= 24'd713764;
        711: data_ff <= -24'd400944;
        712: data_ff <= 24'd222471;
        713: data_ff <= -24'd117134;
        714: data_ff <= 24'd56834;
        715: data_ff <= -24'd24663;
        716: data_ff <= 24'd9203;
        717: data_ff <= -24'd2770;
        718: data_ff <= 24'd581;
        719: data_ff <= -24'd42;
        720: data_ff <= 24'd3929047;
        721: data_ff <= -24'd1381305;
        722: data_ff <= 24'd721951;
        723: data_ff <= -24'd405433;
        724: data_ff <= 24'd224976;
        725: data_ff <= -24'd118484;
        726: data_ff <= 24'd57514;
        727: data_ff <= -24'd24975;
        728: data_ff <= 24'd9328;
        729: data_ff <= -24'd2812;
        730: data_ff <= 24'd592;
        731: data_ff <= -24'd43;
        732: data_ff <= 24'd4000318;
        733: data_ff <= -24'd1398092;
        734: data_ff <= 24'd729911;
        735: data_ff <= -24'd409794;
        736: data_ff <= 24'd227410;
        737: data_ff <= -24'd119798;
        738: data_ff <= 24'd58177;
        739: data_ff <= -24'd25279;
        740: data_ff <= 24'd9451;
        741: data_ff <= -24'd2853;
        742: data_ff <= 24'd602;
        743: data_ff <= -24'd45;
        744: data_ff <= 24'd4071507;
        745: data_ff <= -24'd1414485;
        746: data_ff <= 24'd737642;
        747: data_ff <= -24'd414022;
        748: data_ff <= 24'd229771;
        749: data_ff <= -24'd121073;
        750: data_ff <= 24'd58823;
        751: data_ff <= -24'd25576;
        752: data_ff <= 24'd9571;
        753: data_ff <= -24'd2894;
        754: data_ff <= 24'd613;
        755: data_ff <= -24'd46;
        756: data_ff <= 24'd4142597;
        757: data_ff <= -24'd1430472;
        758: data_ff <= 24'd745138;
        759: data_ff <= -24'd418116;
        760: data_ff <= 24'd232058;
        761: data_ff <= -24'd122311;
        762: data_ff <= 24'd59450;
        763: data_ff <= -24'd25866;
        764: data_ff <= 24'd9688;
        765: data_ff <= -24'd2934;
        766: data_ff <= 24'd623;
        767: data_ff <= -24'd47;
        768: data_ff <= 24'd4213573;
        769: data_ff <= -24'd1446043;
        770: data_ff <= 24'd752394;
        771: data_ff <= -24'd422073;
        772: data_ff <= 24'd234269;
        773: data_ff <= -24'd123509;
        774: data_ff <= 24'd60060;
        775: data_ff <= -24'd26148;
        776: data_ff <= 24'd9803;
        777: data_ff <= -24'd2973;
        778: data_ff <= 24'd633;
        779: data_ff <= -24'd49;
        780: data_ff <= 24'd4284420;
        781: data_ff <= -24'd1461191;
        782: data_ff <= 24'd759407;
        783: data_ff <= -24'd425891;
        784: data_ff <= 24'd236403;
        785: data_ff <= -24'd124668;
        786: data_ff <= 24'd60650;
        787: data_ff <= -24'd26422;
        788: data_ff <= 24'd9915;
        789: data_ff <= -24'd3011;
        790: data_ff <= 24'd643;
        791: data_ff <= -24'd50;
        792: data_ff <= 24'd4355121;
        793: data_ff <= -24'd1475903;
        794: data_ff <= 24'd766170;
        795: data_ff <= -24'd429566;
        796: data_ff <= 24'd238458;
        797: data_ff <= -24'd125785;
        798: data_ff <= 24'd61221;
        799: data_ff <= -24'd26688;
        800: data_ff <= 24'd10025;
        801: data_ff <= -24'd3049;
        802: data_ff <= 24'd653;
        803: data_ff <= -24'd52;
        804: data_ff <= 24'd4425662;
        805: data_ff <= -24'd1490172;
        806: data_ff <= 24'd772680;
        807: data_ff <= -24'd433096;
        808: data_ff <= 24'd240434;
        809: data_ff <= -24'd126861;
        810: data_ff <= 24'd61772;
        811: data_ff <= -24'd26946;
        812: data_ff <= 24'd10131;
        813: data_ff <= -24'd3086;
        814: data_ff <= 24'd663;
        815: data_ff <= -24'd53;
        816: data_ff <= 24'd4496026;
        817: data_ff <= -24'd1503988;
        818: data_ff <= 24'd778933;
        819: data_ff <= -24'd436480;
        820: data_ff <= 24'd242327;
        821: data_ff <= -24'd127895;
        822: data_ff <= 24'd62303;
        823: data_ff <= -24'd27195;
        824: data_ff <= 24'd10234;
        825: data_ff <= -24'd3122;
        826: data_ff <= 24'd673;
        827: data_ff <= -24'd54;
        828: data_ff <= 24'd4566199;
        829: data_ff <= -24'd1517340;
        830: data_ff <= 24'd784923;
        831: data_ff <= -24'd439714;
        832: data_ff <= 24'd244138;
        833: data_ff <= -24'd128885;
        834: data_ff <= 24'd62813;
        835: data_ff <= -24'd27435;
        836: data_ff <= 24'd10334;
        837: data_ff <= -24'd3157;
        838: data_ff <= 24'd682;
        839: data_ff <= -24'd56;
        840: data_ff <= 24'd4636164;
        841: data_ff <= -24'd1530220;
        842: data_ff <= 24'd790647;
        843: data_ff <= -24'd442795;
        844: data_ff <= 24'd245865;
        845: data_ff <= -24'd129831;
        846: data_ff <= 24'd63302;
        847: data_ff <= -24'd27667;
        848: data_ff <= 24'd10431;
        849: data_ff <= -24'd3191;
        850: data_ff <= 24'd692;
        851: data_ff <= -24'd57;
        852: data_ff <= 24'd4705906;
        853: data_ff <= -24'd1542619;
        854: data_ff <= 24'd796101;
        855: data_ff <= -24'd445723;
        856: data_ff <= 24'd247506;
        857: data_ff <= -24'd130733;
        858: data_ff <= 24'd63770;
        859: data_ff <= -24'd27889;
        860: data_ff <= 24'd10525;
        861: data_ff <= -24'd3225;
        862: data_ff <= 24'd701;
        863: data_ff <= -24'd59;
        864: data_ff <= 24'd4775409;
        865: data_ff <= -24'd1554527;
        866: data_ff <= 24'd801280;
        867: data_ff <= -24'd448494;
        868: data_ff <= 24'd249060;
        869: data_ff <= -24'd131589;
        870: data_ff <= 24'd64216;
        871: data_ff <= -24'd28103;
        872: data_ff <= 24'd10616;
        873: data_ff <= -24'd3257;
        874: data_ff <= 24'd710;
        875: data_ff <= -24'd60;
        876: data_ff <= 24'd4844659;
        877: data_ff <= -24'd1565934;
        878: data_ff <= 24'd806180;
        879: data_ff <= -24'd451107;
        880: data_ff <= 24'd250526;
        881: data_ff <= -24'd132399;
        882: data_ff <= 24'd64640;
        883: data_ff <= -24'd28306;
        884: data_ff <= 24'd10702;
        885: data_ff <= -24'd3288;
        886: data_ff <= 24'd719;
        887: data_ff <= -24'd62;
        888: data_ff <= 24'd4913639;
        889: data_ff <= -24'd1576833;
        890: data_ff <= 24'd810797;
        891: data_ff <= -24'd453558;
        892: data_ff <= 24'd251902;
        893: data_ff <= -24'd133161;
        894: data_ff <= 24'd65041;
        895: data_ff <= -24'd28500;
        896: data_ff <= 24'd10786;
        897: data_ff <= -24'd3319;
        898: data_ff <= 24'd728;
        899: data_ff <= -24'd63;
        900: data_ff <= 24'd4982333;
        901: data_ff <= -24'd1587214;
        902: data_ff <= 24'd815127;
        903: data_ff <= -24'd455847;
        904: data_ff <= 24'd253188;
        905: data_ff <= -24'd133877;
        906: data_ff <= 24'd65419;
        907: data_ff <= -24'd28685;
        908: data_ff <= 24'd10866;
        909: data_ff <= -24'd3348;
        910: data_ff <= 24'd736;
        911: data_ff <= -24'd65;
        912: data_ff <= 24'd5050727;
        913: data_ff <= -24'd1597069;
        914: data_ff <= 24'd819167;
        915: data_ff <= -24'd457970;
        916: data_ff <= 24'd254382;
        917: data_ff <= -24'd134544;
        918: data_ff <= 24'd65774;
        919: data_ff <= -24'd28859;
        920: data_ff <= 24'd10942;
        921: data_ff <= -24'd3376;
        922: data_ff <= 24'd745;
        923: data_ff <= -24'd66;
        924: data_ff <= 24'd5118806;
        925: data_ff <= -24'd1606387;
        926: data_ff <= 24'd822912;
        927: data_ff <= -24'd459926;
        928: data_ff <= 24'd255483;
        929: data_ff <= -24'd135161;
        930: data_ff <= 24'd66105;
        931: data_ff <= -24'd29022;
        932: data_ff <= 24'd11014;
        933: data_ff <= -24'd3403;
        934: data_ff <= 24'd753;
        935: data_ff <= -24'd67;
        936: data_ff <= 24'd5186552;
        937: data_ff <= -24'd1615162;
        938: data_ff <= 24'd826360;
        939: data_ff <= -24'd461713;
        940: data_ff <= 24'd256489;
        941: data_ff <= -24'd135729;
        942: data_ff <= 24'd66412;
        943: data_ff <= -24'd29176;
        944: data_ff <= 24'd11082;
        945: data_ff <= -24'd3429;
        946: data_ff <= 24'd760;
        947: data_ff <= -24'd69;
        948: data_ff <= 24'd5253953;
        949: data_ff <= -24'd1623383;
        950: data_ff <= 24'd829505;
        951: data_ff <= -24'd463329;
        952: data_ff <= 24'd257400;
        953: data_ff <= -24'd136247;
        954: data_ff <= 24'd66694;
        955: data_ff <= -24'd29319;
        956: data_ff <= 24'd11147;
        957: data_ff <= -24'd3454;
        958: data_ff <= 24'd768;
        959: data_ff <= -24'd70;
        960: data_ff <= 24'd5320991;
        961: data_ff <= -24'd1631044;
        962: data_ff <= 24'd832346;
        963: data_ff <= -24'd464772;
        964: data_ff <= 24'd258215;
        965: data_ff <= -24'd136714;
        966: data_ff <= 24'd66952;
        967: data_ff <= -24'd29451;
        968: data_ff <= 24'd11207;
        969: data_ff <= -24'd3478;
        970: data_ff <= 24'd775;
        971: data_ff <= -24'd72;
        972: data_ff <= 24'd5387652;
        973: data_ff <= -24'd1638134;
        974: data_ff <= 24'd834878;
        975: data_ff <= -24'd466040;
        976: data_ff <= 24'd258932;
        977: data_ff <= -24'd137129;
        978: data_ff <= 24'd67185;
        979: data_ff <= -24'd29572;
        980: data_ff <= 24'd11264;
        981: data_ff <= -24'd3500;
        982: data_ff <= 24'd783;
        983: data_ff <= -24'd73;
        984: data_ff <= 24'd5453920;
        985: data_ff <= -24'd1644647;
        986: data_ff <= 24'd837098;
        987: data_ff <= -24'd467131;
        988: data_ff <= 24'd259551;
        989: data_ff <= -24'd137492;
        990: data_ff <= 24'd67392;
        991: data_ff <= -24'd29681;
        992: data_ff <= 24'd11316;
        993: data_ff <= -24'd3521;
        994: data_ff <= 24'd789;
        995: data_ff <= -24'd75;
        996: data_ff <= 24'd5519781;
        997: data_ff <= -24'd1650574;
        998: data_ff <= 24'd839004;
        999: data_ff <= -24'd468045;
        1000: data_ff <= 24'd260070;
        1001: data_ff <= -24'd137803;
        1002: data_ff <= 24'd67573;
        1003: data_ff <= -24'd29780;
        1004: data_ff <= 24'd11364;
        1005: data_ff <= -24'd3541;
        1006: data_ff <= 24'd796;
        1007: data_ff <= -24'd76;
        1008: data_ff <= 24'd5585220;
        1009: data_ff <= -24'd1655907;
        1010: data_ff <= 24'd840590;
        1011: data_ff <= -24'd468778;
        1012: data_ff <= 24'd260489;
        1013: data_ff <= -24'd138060;
        1014: data_ff <= 24'd67728;
        1015: data_ff <= -24'd29867;
        1016: data_ff <= 24'd11407;
        1017: data_ff <= -24'd3560;
        1018: data_ff <= 24'd802;
        1019: data_ff <= -24'd77;
        1020: data_ff <= 24'd5650221;
        1021: data_ff <= -24'd1660638;
        1022: data_ff <= 24'd841856;
        1023: data_ff <= -24'd469330;
        1024: data_ff <= 24'd260807;
        1025: data_ff <= -24'd138263;
        1026: data_ff <= 24'd67857;
        1027: data_ff <= -24'd29943;
        1028: data_ff <= 24'd11446;
        1029: data_ff <= -24'd3577;
        1030: data_ff <= 24'd808;
        1031: data_ff <= -24'd79;
        1032: data_ff <= 24'd5714769;
        1033: data_ff <= -24'd1664760;
        1034: data_ff <= 24'd842798;
        1035: data_ff <= -24'd469699;
        1036: data_ff <= 24'd261022;
        1037: data_ff <= -24'd138411;
        1038: data_ff <= 24'd67959;
        1039: data_ff <= -24'd30006;
        1040: data_ff <= 24'd11481;
        1041: data_ff <= -24'd3593;
        1042: data_ff <= 24'd814;
        1043: data_ff <= -24'd80;
        1044: data_ff <= 24'd5778850;
        1045: data_ff <= -24'd1668264;
        1046: data_ff <= 24'd843412;
        1047: data_ff <= -24'd469883;
        1048: data_ff <= 24'd261134;
        1049: data_ff <= -24'd138505;
        1050: data_ff <= 24'd68033;
        1051: data_ff <= -24'd30058;
        1052: data_ff <= 24'd11511;
        1053: data_ff <= -24'd3607;
        1054: data_ff <= 24'd819;
        1055: data_ff <= -24'd81;
        1056: data_ff <= 24'd5842449;
        1057: data_ff <= -24'd1671144;
        1058: data_ff <= 24'd843697;
        1059: data_ff <= -24'd469882;
        1060: data_ff <= 24'd261142;
        1061: data_ff <= -24'd138543;
        1062: data_ff <= 24'd68081;
        1063: data_ff <= -24'd30097;
        1064: data_ff <= 24'd11537;
        1065: data_ff <= -24'd3620;
        1066: data_ff <= 24'd824;
        1067: data_ff <= -24'd83;
        1068: data_ff <= 24'd5905552;
        1069: data_ff <= -24'd1673392;
        1070: data_ff <= 24'd843650;
        1071: data_ff <= -24'd469694;
        1072: data_ff <= 24'd261045;
        1073: data_ff <= -24'd138526;
        1074: data_ff <= 24'd68101;
        1075: data_ff <= -24'd30125;
        1076: data_ff <= 24'd11557;
        1077: data_ff <= -24'd3632;
        1078: data_ff <= 24'd829;
        1079: data_ff <= -24'd84;
        1080: data_ff <= 24'd5968143;
        1081: data_ff <= -24'd1675000;
        1082: data_ff <= 24'd843268;
        1083: data_ff <= -24'd469317;
        1084: data_ff <= 24'd260843;
        1085: data_ff <= -24'd138452;
        1086: data_ff <= 24'd68093;
        1087: data_ff <= -24'd30140;
        1088: data_ff <= 24'd11573;
        1089: data_ff <= -24'd3642;
        1090: data_ff <= 24'd834;
        1091: data_ff <= -24'd85;
        1092: data_ff <= 24'd6030208;
        1093: data_ff <= -24'd1675962;
        1094: data_ff <= 24'd842548;
        1095: data_ff <= -24'd468750;
        1096: data_ff <= 24'd260534;
        1097: data_ff <= -24'd138321;
        1098: data_ff <= 24'd68057;
        1099: data_ff <= -24'd30142;
        1100: data_ff <= 24'd11585;
        1101: data_ff <= -24'd3650;
        1102: data_ff <= 24'd838;
        1103: data_ff <= -24'd87;
        1104: data_ff <= 24'd6091733;
        1105: data_ff <= -24'd1676270;
        1106: data_ff <= 24'd841489;
        1107: data_ff <= -24'd467993;
        1108: data_ff <= 24'd260119;
        1109: data_ff <= -24'd138133;
        1110: data_ff <= 24'd67992;
        1111: data_ff <= -24'd30132;
        1112: data_ff <= 24'd11591;
        1113: data_ff <= -24'd3657;
        1114: data_ff <= 24'd841;
        1115: data_ff <= -24'd88;
        1116: data_ff <= 24'd6152704;
        1117: data_ff <= -24'd1675918;
        1118: data_ff <= 24'd840089;
        1119: data_ff <= -24'd467043;
        1120: data_ff <= 24'd259596;
        1121: data_ff <= -24'd137888;
        1122: data_ff <= 24'd67899;
        1123: data_ff <= -24'd30109;
        1124: data_ff <= 24'd11592;
        1125: data_ff <= -24'd3662;
        1126: data_ff <= 24'd845;
        1127: data_ff <= -24'd89;
        1128: data_ff <= 24'd6213106;
        1129: data_ff <= -24'd1674900;
        1130: data_ff <= 24'd838344;
        1131: data_ff <= -24'd465901;
        1132: data_ff <= 24'd258965;
        1133: data_ff <= -24'd137584;
        1134: data_ff <= 24'd67777;
        1135: data_ff <= -24'd30073;
        1136: data_ff <= 24'd11588;
        1137: data_ff <= -24'd3666;
        1138: data_ff <= 24'd848;
        1139: data_ff <= -24'd90;
        1140: data_ff <= 24'd6272925;
        1141: data_ff <= -24'd1673208;
        1142: data_ff <= 24'd836255;
        1143: data_ff <= -24'd464565;
        1144: data_ff <= 24'd258225;
        1145: data_ff <= -24'd137222;
        1146: data_ff <= 24'd67626;
        1147: data_ff <= -24'd30023;
        1148: data_ff <= 24'd11579;
        1149: data_ff <= -24'd3668;
        1150: data_ff <= 24'd850;
        1151: data_ff <= -24'd91;
        1152: data_ff <= 24'd6332148;
        1153: data_ff <= -24'd1670836;
        1154: data_ff <= 24'd833817;
        1155: data_ff <= -24'd463035;
        1156: data_ff <= 24'd257376;
        1157: data_ff <= -24'd136802;
        1158: data_ff <= 24'd67446;
        1159: data_ff <= -24'd29961;
        1160: data_ff <= 24'd11565;
        1161: data_ff <= -24'd3668;
        1162: data_ff <= 24'd852;
        1163: data_ff <= -24'd92;
        1164: data_ff <= 24'd6390760;
        1165: data_ff <= -24'd1667779;
        1166: data_ff <= 24'd831030;
        1167: data_ff <= -24'd461309;
        1168: data_ff <= 24'd256418;
        1169: data_ff <= -24'd136322;
        1170: data_ff <= 24'd67236;
        1171: data_ff <= -24'd29886;
        1172: data_ff <= 24'd11546;
        1173: data_ff <= -24'd3667;
        1174: data_ff <= 24'd854;
        1175: data_ff <= -24'd93;
        1176: data_ff <= 24'd6448748;
        1177: data_ff <= -24'd1664030;
        1178: data_ff <= 24'd827893;
        1179: data_ff <= -24'd459386;
        1180: data_ff <= 24'd255349;
        1181: data_ff <= -24'd135784;
        1182: data_ff <= 24'd66996;
        1183: data_ff <= -24'd29796;
        1184: data_ff <= 24'd11521;
        1185: data_ff <= -24'd3664;
        1186: data_ff <= 24'd856;
        1187: data_ff <= -24'd94;
        1188: data_ff <= 24'd6506099;
        1189: data_ff <= -24'd1659583;
        1190: data_ff <= 24'd824403;
        1191: data_ff <= -24'd457268;
        1192: data_ff <= 24'd254170;
        1193: data_ff <= -24'd135185;
        1194: data_ff <= 24'd66727;
        1195: data_ff <= -24'd29694;
        1196: data_ff <= 24'd11492;
        1197: data_ff <= -24'd3659;
        1198: data_ff <= 24'd857;
        1199: data_ff <= -24'd95;
        1200: data_ff <= 24'd6562798;
        1201: data_ff <= -24'd1654433;
        1202: data_ff <= 24'd820560;
        1203: data_ff <= -24'd454951;
        1204: data_ff <= 24'd252880;
        1205: data_ff <= -24'd134527;
        1206: data_ff <= 24'd66428;
        1207: data_ff <= -24'd29578;
        1208: data_ff <= 24'd11456;
        1209: data_ff <= -24'd3653;
        1210: data_ff <= 24'd857;
        1211: data_ff <= -24'd96;
        1212: data_ff <= 24'd6618833;
        1213: data_ff <= -24'd1648573;
        1214: data_ff <= 24'd816362;
        1215: data_ff <= -24'd452437;
        1216: data_ff <= 24'd251479;
        1217: data_ff <= -24'd133809;
        1218: data_ff <= 24'd66098;
        1219: data_ff <= -24'd29448;
        1220: data_ff <= 24'd11415;
        1221: data_ff <= -24'd3644;
        1222: data_ff <= 24'd857;
        1223: data_ff <= -24'd97;
        1224: data_ff <= 24'd6674190;
        1225: data_ff <= -24'd1642000;
        1226: data_ff <= 24'd811808;
        1227: data_ff <= -24'd449725;
        1228: data_ff <= 24'd249967;
        1229: data_ff <= -24'd133031;
        1230: data_ff <= 24'd65738;
        1231: data_ff <= -24'd29304;
        1232: data_ff <= 24'd11369;
        1233: data_ff <= -24'd3634;
        1234: data_ff <= 24'd857;
        1235: data_ff <= -24'd97;
        1236: data_ff <= 24'd6728856;
        1237: data_ff <= -24'd1634707;
        1238: data_ff <= 24'd806897;
        1239: data_ff <= -24'd446813;
        1240: data_ff <= 24'd248343;
        1241: data_ff <= -24'd132192;
        1242: data_ff <= 24'd65348;
        1243: data_ff <= -24'd29147;
        1244: data_ff <= 24'd11317;
        1245: data_ff <= -24'd3622;
        1246: data_ff <= 24'd856;
        1247: data_ff <= -24'd98;
        1248: data_ff <= 24'd6782819;
        1249: data_ff <= -24'd1626689;
        1250: data_ff <= 24'd801629;
        1251: data_ff <= -24'd443703;
        1252: data_ff <= 24'd246607;
        1253: data_ff <= -24'd131293;
        1254: data_ff <= 24'd64927;
        1255: data_ff <= -24'd28975;
        1256: data_ff <= 24'd11260;
        1257: data_ff <= -24'd3609;
        1258: data_ff <= 24'd855;
        1259: data_ff <= -24'd99;
        1260: data_ff <= 24'd6836066;
        1261: data_ff <= -24'd1617942;
        1262: data_ff <= 24'd796002;
        1263: data_ff <= -24'd440394;
        1264: data_ff <= 24'd244759;
        1265: data_ff <= -24'd130334;
        1266: data_ff <= 24'd64476;
        1267: data_ff <= -24'd28789;
        1268: data_ff <= 24'd11197;
        1269: data_ff <= -24'd3593;
        1270: data_ff <= 24'd853;
        1271: data_ff <= -24'd99;
        1272: data_ff <= 24'd6888584;
        1273: data_ff <= -24'd1608461;
        1274: data_ff <= 24'd790016;
        1275: data_ff <= -24'd436886;
        1276: data_ff <= 24'd242799;
        1277: data_ff <= -24'd129313;
        1278: data_ff <= 24'd63994;
        1279: data_ff <= -24'd28590;
        1280: data_ff <= 24'd11128;
        1281: data_ff <= -24'd3575;
        1282: data_ff <= 24'd851;
        1283: data_ff <= -24'd100;
        1284: data_ff <= 24'd6940360;
        1285: data_ff <= -24'd1598241;
        1286: data_ff <= 24'd783670;
        1287: data_ff <= -24'd433179;
        1288: data_ff <= 24'd240727;
        1289: data_ff <= -24'd128232;
        1290: data_ff <= 24'd63481;
        1291: data_ff <= -24'd28376;
        1292: data_ff <= 24'd11054;
        1293: data_ff <= -24'd3556;
        1294: data_ff <= 24'd848;
        1295: data_ff <= -24'd100;
        1296: data_ff <= 24'd6991383;
        1297: data_ff <= -24'd1587279;
        1298: data_ff <= 24'd776965;
        1299: data_ff <= -24'd429272;
        1300: data_ff <= 24'd238543;
        1301: data_ff <= -24'd127090;
        1302: data_ff <= 24'd62937;
        1303: data_ff <= -24'd28148;
        1304: data_ff <= 24'd10974;
        1305: data_ff <= -24'd3534;
        1306: data_ff <= 24'd845;
        1307: data_ff <= -24'd101;
        1308: data_ff <= 24'd7041641;
        1309: data_ff <= -24'd1575569;
        1310: data_ff <= 24'd769900;
        1311: data_ff <= -24'd425166;
        1312: data_ff <= 24'd236247;
        1313: data_ff <= -24'd125887;
        1314: data_ff <= 24'd62362;
        1315: data_ff <= -24'd27905;
        1316: data_ff <= 24'd10888;
        1317: data_ff <= -24'd3511;
        1318: data_ff <= 24'd841;
        1319: data_ff <= -24'd101;
        1320: data_ff <= 24'd7091121;
        1321: data_ff <= -24'd1563109;
        1322: data_ff <= 24'd762475;
        1323: data_ff <= -24'd420862;
        1324: data_ff <= 24'd233839;
        1325: data_ff <= -24'd124623;
        1326: data_ff <= 24'd61756;
        1327: data_ff <= -24'd27648;
        1328: data_ff <= 24'd10796;
        1329: data_ff <= -24'd3485;
        1330: data_ff <= 24'd837;
        1331: data_ff <= -24'd101;
        1332: data_ff <= 24'd7139811;
        1333: data_ff <= -24'd1549894;
        1334: data_ff <= 24'd754690;
        1335: data_ff <= -24'd416359;
        1336: data_ff <= 24'd231319;
        1337: data_ff <= -24'd123298;
        1338: data_ff <= 24'd61119;
        1339: data_ff <= -24'd27377;
        1340: data_ff <= 24'd10698;
        1341: data_ff <= -24'd3458;
        1342: data_ff <= 24'd832;
        1343: data_ff <= -24'd102;
        1344: data_ff <= 24'd7187701;
        1345: data_ff <= -24'd1535921;
        1346: data_ff <= 24'd746545;
        1347: data_ff <= -24'd411657;
        1348: data_ff <= 24'd228688;
        1349: data_ff <= -24'd121912;
        1350: data_ff <= 24'd60451;
        1351: data_ff <= -24'd27092;
        1352: data_ff <= 24'd10595;
        1353: data_ff <= -24'd3429;
        1354: data_ff <= 24'd827;
        1355: data_ff <= -24'd102;
        1356: data_ff <= 24'd7234779;
        1357: data_ff <= -24'd1521187;
        1358: data_ff <= 24'd738041;
        1359: data_ff <= -24'd406758;
        1360: data_ff <= 24'd225945;
        1361: data_ff <= -24'd120466;
        1362: data_ff <= 24'd59752;
        1363: data_ff <= -24'd26791;
        1364: data_ff <= 24'd10485;
        1365: data_ff <= -24'd3397;
        1366: data_ff <= 24'd821;
        1367: data_ff <= -24'd102;
        1368: data_ff <= 24'd7281033;
        1369: data_ff <= -24'd1505688;
        1370: data_ff <= 24'd729179;
        1371: data_ff <= -24'd401662;
        1372: data_ff <= 24'd223091;
        1373: data_ff <= -24'd118958;
        1374: data_ff <= 24'd59022;
        1375: data_ff <= -24'd26477;
        1376: data_ff <= 24'd10370;
        1377: data_ff <= -24'd3364;
        1378: data_ff <= 24'd815;
        1379: data_ff <= -24'd102;
        1380: data_ff <= 24'd7326453;
        1381: data_ff <= -24'd1489422;
        1382: data_ff <= 24'd719958;
        1383: data_ff <= -24'd396369;
        1384: data_ff <= 24'd220126;
        1385: data_ff <= -24'd117391;
        1386: data_ff <= 24'd58261;
        1387: data_ff <= -24'd26148;
        1388: data_ff <= 24'd10248;
        1389: data_ff <= -24'd3328;
        1390: data_ff <= 24'd808;
        1391: data_ff <= -24'd101;
        1392: data_ff <= 24'd7371027;
        1393: data_ff <= -24'd1472385;
        1394: data_ff <= 24'd710380;
        1395: data_ff <= -24'd390880;
        1396: data_ff <= 24'd217051;
        1397: data_ff <= -24'd115763;
        1398: data_ff <= 24'd57469;
        1399: data_ff <= -24'd25804;
        1400: data_ff <= 24'd10121;
        1401: data_ff <= -24'd3290;
        1402: data_ff <= 24'd801;
        1403: data_ff <= -24'd101;
        1404: data_ff <= 24'd7414746;
        1405: data_ff <= -24'd1454575;
        1406: data_ff <= 24'd700445;
        1407: data_ff <= -24'd385196;
        1408: data_ff <= 24'd213866;
        1409: data_ff <= -24'd114074;
        1410: data_ff <= 24'd56646;
        1411: data_ff <= -24'd25446;
        1412: data_ff <= 24'd9987;
        1413: data_ff <= -24'd3251;
        1414: data_ff <= 24'd793;
        1415: data_ff <= -24'd101;
        1416: data_ff <= 24'd7457598;
        1417: data_ff <= -24'd1435990;
        1418: data_ff <= 24'd690155;
        1419: data_ff <= -24'd379318;
        1420: data_ff <= 24'd210572;
        1421: data_ff <= -24'd112326;
        1422: data_ff <= 24'd55792;
        1423: data_ff <= -24'd25073;
        1424: data_ff <= 24'd9848;
        1425: data_ff <= -24'd3209;
        1426: data_ff <= 24'd784;
        1427: data_ff <= -24'd101;
        1428: data_ff <= 24'd7499573;
        1429: data_ff <= -24'd1416628;
        1430: data_ff <= 24'd679511;
        1431: data_ff <= -24'd373246;
        1432: data_ff <= 24'd207169;
        1433: data_ff <= -24'd110518;
        1434: data_ff <= 24'd54907;
        1435: data_ff <= -24'd24686;
        1436: data_ff <= 24'd9702;
        1437: data_ff <= -24'd3165;
        1438: data_ff <= 24'd775;
        1439: data_ff <= -24'd100;
        1440: data_ff <= 24'd7540662;
        1441: data_ff <= -24'd1396487;
        1442: data_ff <= 24'd668514;
        1443: data_ff <= -24'd366982;
        1444: data_ff <= 24'd203657;
        1445: data_ff <= -24'd108650;
        1446: data_ff <= 24'd53991;
        1447: data_ff <= -24'd24285;
        1448: data_ff <= 24'd9551;
        1449: data_ff <= -24'd3119;
        1450: data_ff <= 24'd765;
        1451: data_ff <= -24'd99;
        1452: data_ff <= 24'd7580855;
        1453: data_ff <= -24'd1375564;
        1454: data_ff <= 24'd657165;
        1455: data_ff <= -24'd360527;
        1456: data_ff <= 24'd200037;
        1457: data_ff <= -24'd106723;
        1458: data_ff <= 24'd53045;
        1459: data_ff <= -24'd23868;
        1460: data_ff <= 24'd9393;
        1461: data_ff <= -24'd3070;
        1462: data_ff <= 24'd755;
        1463: data_ff <= -24'd99;
        1464: data_ff <= 24'd7620141;
        1465: data_ff <= -24'd1353859;
        1466: data_ff <= 24'd645467;
        1467: data_ff <= -24'd353882;
        1468: data_ff <= 24'd196310;
        1469: data_ff <= -24'd104738;
        1470: data_ff <= 24'd52068;
        1471: data_ff <= -24'd23438;
        1472: data_ff <= 24'd9229;
        1473: data_ff <= -24'd3020;
        1474: data_ff <= 24'd744;
        1475: data_ff <= -24'd98;
        1476: data_ff <= 24'd7658511;
        1477: data_ff <= -24'd1331371;
        1478: data_ff <= 24'd633422;
        1479: data_ff <= -24'd347048;
        1480: data_ff <= 24'd192477;
        1481: data_ff <= -24'd102693;
        1482: data_ff <= 24'd51061;
        1483: data_ff <= -24'd22993;
        1484: data_ff <= 24'd9060;
        1485: data_ff <= -24'd2968;
        1486: data_ff <= 24'd732;
        1487: data_ff <= -24'd97;
        1488: data_ff <= 24'd7695957;
        1489: data_ff <= -24'd1308097;
        1490: data_ff <= 24'd621030;
        1491: data_ff <= -24'd340027;
        1492: data_ff <= 24'd188538;
        1493: data_ff <= -24'd100591;
        1494: data_ff <= 24'd50024;
        1495: data_ff <= -24'd22533;
        1496: data_ff <= 24'd8884;
        1497: data_ff <= -24'd2913;
        1498: data_ff <= 24'd720;
        1499: data_ff <= -24'd96;
        1500: data_ff <= 24'd7732469;
        1501: data_ff <= -24'd1284038;
        1502: data_ff <= 24'd608294;
        1503: data_ff <= -24'd332819;
        1504: data_ff <= 24'd184494;
        1505: data_ff <= -24'd98430;
        1506: data_ff <= 24'd48956;
        1507: data_ff <= -24'd22060;
        1508: data_ff <= 24'd8702;
        1509: data_ff <= -24'd2856;
        1510: data_ff <= 24'd707;
        1511: data_ff <= -24'd95;
        1512: data_ff <= 24'd7768038;
        1513: data_ff <= -24'd1259192;
        1514: data_ff <= 24'd595216;
        1515: data_ff <= -24'd325427;
        1516: data_ff <= 24'd180346;
        1517: data_ff <= -24'd96212;
        1518: data_ff <= 24'd47859;
        1519: data_ff <= -24'd21572;
        1520: data_ff <= 24'd8514;
        1521: data_ff <= -24'd2797;
        1522: data_ff <= 24'd694;
        1523: data_ff <= -24'd94;
        1524: data_ff <= 24'd7802657;
        1525: data_ff <= -24'd1233560;
        1526: data_ff <= 24'd581799;
        1527: data_ff <= -24'd317853;
        1528: data_ff <= 24'd176095;
        1529: data_ff <= -24'd93937;
        1530: data_ff <= 24'd46732;
        1531: data_ff <= -24'd21069;
        1532: data_ff <= 24'd8320;
        1533: data_ff <= -24'd2736;
        1534: data_ff <= 24'd680;
        1535: data_ff <= -24'd92;
        1536: data_ff <= 24'd7836316;
        1537: data_ff <= -24'd1207140;
        1538: data_ff <= 24'd568046;
        1539: data_ff <= -24'd310097;
        1540: data_ff <= 24'd171742;
        1541: data_ff <= -24'd91606;
        1542: data_ff <= 24'd45575;
        1543: data_ff <= -24'd20553;
        1544: data_ff <= 24'd8120;
        1545: data_ff <= -24'd2672;
        1546: data_ff <= 24'd665;
        1547: data_ff <= -24'd91;
        1548: data_ff <= 24'd7869007;
        1549: data_ff <= -24'd1179934;
        1550: data_ff <= 24'd553958;
        1551: data_ff <= -24'd302162;
        1552: data_ff <= 24'd167288;
        1553: data_ff <= -24'd89219;
        1554: data_ff <= 24'd44389;
        1555: data_ff <= -24'd20022;
        1556: data_ff <= 24'd7914;
        1557: data_ff <= -24'd2607;
        1558: data_ff <= 24'd650;
        1559: data_ff <= -24'd89;
        1560: data_ff <= 24'd7900723;
        1561: data_ff <= -24'd1151940;
        1562: data_ff <= 24'd539538;
        1563: data_ff <= -24'd294049;
        1564: data_ff <= 24'd162734;
        1565: data_ff <= -24'd86776;
        1566: data_ff <= 24'd43174;
        1567: data_ff <= -24'd19478;
        1568: data_ff <= 24'd7702;
        1569: data_ff <= -24'd2539;
        1570: data_ff <= 24'd634;
        1571: data_ff <= -24'd88;
        1572: data_ff <= 24'd7931455;
        1573: data_ff <= -24'd1123160;
        1574: data_ff <= 24'd524790;
        1575: data_ff <= -24'd285761;
        1576: data_ff <= 24'd158080;
        1577: data_ff <= -24'd84278;
        1578: data_ff <= 24'd41930;
        1579: data_ff <= -24'd18919;
        1580: data_ff <= 24'd7484;
        1581: data_ff <= -24'd2469;
        1582: data_ff <= 24'd618;
        1583: data_ff <= -24'd86;
        1584: data_ff <= 24'd7961198;
        1585: data_ff <= -24'd1093594;
        1586: data_ff <= 24'd509717;
        1587: data_ff <= -24'd277299;
        1588: data_ff <= 24'd153329;
        1589: data_ff <= -24'd81726;
        1590: data_ff <= 24'd40657;
        1591: data_ff <= -24'd18347;
        1592: data_ff <= 24'd7260;
        1593: data_ff <= -24'd2397;
        1594: data_ff <= 24'd601;
        1595: data_ff <= -24'd84;
        1596: data_ff <= 24'd7989942;
        1597: data_ff <= -24'd1063244;
        1598: data_ff <= 24'd494322;
        1599: data_ff <= -24'd268666;
        1600: data_ff <= 24'd148481;
        1601: data_ff <= -24'd79120;
        1602: data_ff <= 24'd39356;
        1603: data_ff <= -24'd17761;
        1604: data_ff <= 24'd7030;
        1605: data_ff <= -24'd2322;
        1606: data_ff <= 24'd583;
        1607: data_ff <= -24'd82;
        1608: data_ff <= 24'd8017682;
        1609: data_ff <= -24'd1032109;
        1610: data_ff <= 24'd478608;
        1611: data_ff <= -24'd259863;
        1612: data_ff <= 24'd143537;
        1613: data_ff <= -24'd76461;
        1614: data_ff <= 24'd38027;
        1615: data_ff <= -24'd17161;
        1616: data_ff <= 24'd6794;
        1617: data_ff <= -24'd2246;
        1618: data_ff <= 24'd565;
        1619: data_ff <= -24'd80;
        1620: data_ff <= 24'd8044411;
        1621: data_ff <= -24'd1000193;
        1622: data_ff <= 24'd462578;
        1623: data_ff <= -24'd250894;
        1624: data_ff <= 24'd138500;
        1625: data_ff <= -24'd73749;
        1626: data_ff <= 24'd36671;
        1627: data_ff <= -24'd16548;
        1628: data_ff <= 24'd6552;
        1629: data_ff <= -24'd2167;
        1630: data_ff <= 24'd546;
        1631: data_ff <= -24'd77;
        1632: data_ff <= 24'd8070121;
        1633: data_ff <= -24'd967495;
        1634: data_ff <= 24'd446237;
        1635: data_ff <= -24'd241760;
        1636: data_ff <= 24'd133370;
        1637: data_ff <= -24'd70986;
        1638: data_ff <= 24'd35287;
        1639: data_ff <= -24'd15921;
        1640: data_ff <= 24'd6305;
        1641: data_ff <= -24'd2086;
        1642: data_ff <= 24'd526;
        1643: data_ff <= -24'd75;
        1644: data_ff <= 24'd8094808;
        1645: data_ff <= -24'd934018;
        1646: data_ff <= 24'd429588;
        1647: data_ff <= -24'd232464;
        1648: data_ff <= 24'd128148;
        1649: data_ff <= -24'd68172;
        1650: data_ff <= 24'd33876;
        1651: data_ff <= -24'd15281;
        1652: data_ff <= 24'd6052;
        1653: data_ff <= -24'd2003;
        1654: data_ff <= 24'd505;
        1655: data_ff <= -24'd72;
        1656: data_ff <= 24'd8118465;
        1657: data_ff <= -24'd899764;
        1658: data_ff <= 24'd412636;
        1659: data_ff <= -24'd223008;
        1660: data_ff <= 24'd122836;
        1661: data_ff <= -24'd65307;
        1662: data_ff <= 24'd32438;
        1663: data_ff <= -24'd14628;
        1664: data_ff <= 24'd5792;
        1665: data_ff <= -24'd1918;
        1666: data_ff <= 24'd484;
        1667: data_ff <= -24'd70;
        1668: data_ff <= 24'd8141086;
        1669: data_ff <= -24'd864735;
        1670: data_ff <= 24'd395383;
        1671: data_ff <= -24'd213395;
        1672: data_ff <= 24'd117436;
        1673: data_ff <= -24'd62393;
        1674: data_ff <= 24'd30973;
        1675: data_ff <= -24'd13963;
        1676: data_ff <= 24'd5528;
        1677: data_ff <= -24'd1830;
        1678: data_ff <= 24'd463;
        1679: data_ff <= -24'd67;
        1680: data_ff <= 24'd8162666;
        1681: data_ff <= -24'd828933;
        1682: data_ff <= 24'd377836;
        1683: data_ff <= -24'd203627;
        1684: data_ff <= 24'd111948;
        1685: data_ff <= -24'd59431;
        1686: data_ff <= 24'd29483;
        1687: data_ff <= -24'd13284;
        1688: data_ff <= 24'd5257;
        1689: data_ff <= -24'd1741;
        1690: data_ff <= 24'd440;
        1691: data_ff <= -24'd64;
        1692: data_ff <= 24'd8183199;
        1693: data_ff <= -24'd792362;
        1694: data_ff <= 24'd359997;
        1695: data_ff <= -24'd193709;
        1696: data_ff <= 24'd106376;
        1697: data_ff <= -24'd56420;
        1698: data_ff <= 24'd27967;
        1699: data_ff <= -24'd12592;
        1700: data_ff <= 24'd4981;
        1701: data_ff <= -24'd1649;
        1702: data_ff <= 24'd418;
        1703: data_ff <= -24'd61;
        1704: data_ff <= 24'd8202681;
        1705: data_ff <= -24'd755023;
        1706: data_ff <= 24'd341871;
        1707: data_ff <= -24'd183641;
        1708: data_ff <= 24'd100719;
        1709: data_ff <= -24'd53362;
        1710: data_ff <= 24'd26426;
        1711: data_ff <= -24'd11888;
        1712: data_ff <= 24'd4699;
        1713: data_ff <= -24'd1555;
        1714: data_ff <= 24'd394;
        1715: data_ff <= -24'd58;
        1716: data_ff <= 24'd8221107;
        1717: data_ff <= -24'd716921;
        1718: data_ff <= 24'd323463;
        1719: data_ff <= -24'd173427;
        1720: data_ff <= 24'd94981;
        1721: data_ff <= -24'd50258;
        1722: data_ff <= 24'd24860;
        1723: data_ff <= -24'd11172;
        1724: data_ff <= 24'd4412;
        1725: data_ff <= -24'd1459;
        1726: data_ff <= 24'd370;
        1727: data_ff <= -24'd54;
        1728: data_ff <= 24'd8238473;
        1729: data_ff <= -24'd678059;
        1730: data_ff <= 24'd304779;
        1731: data_ff <= -24'd163071;
        1732: data_ff <= 24'd89161;
        1733: data_ff <= -24'd47109;
        1734: data_ff <= 24'd23269;
        1735: data_ff <= -24'd10443;
        1736: data_ff <= 24'd4120;
        1737: data_ff <= -24'd1361;
        1738: data_ff <= 24'd345;
        1739: data_ff <= -24'd51;
        1740: data_ff <= 24'd8254773;
        1741: data_ff <= -24'd638439;
        1742: data_ff <= 24'd285822;
        1743: data_ff <= -24'd152574;
        1744: data_ff <= 24'd83264;
        1745: data_ff <= -24'd43915;
        1746: data_ff <= 24'd21655;
        1747: data_ff <= -24'd9703;
        1748: data_ff <= 24'd3822;
        1749: data_ff <= -24'd1261;
        1750: data_ff <= 24'd319;
        1751: data_ff <= -24'd47;
        1752: data_ff <= 24'd8270005;
        1753: data_ff <= -24'd598067;
        1754: data_ff <= 24'd266598;
        1755: data_ff <= -24'd141941;
        1756: data_ff <= 24'd77289;
        1757: data_ff <= -24'd40678;
        1758: data_ff <= 24'd20017;
        1759: data_ff <= -24'd8951;
        1760: data_ff <= 24'd3518;
        1761: data_ff <= -24'd1159;
        1762: data_ff <= 24'd293;
        1763: data_ff <= -24'd43;
        1764: data_ff <= 24'd8284164;
        1765: data_ff <= -24'd556945;
        1766: data_ff <= 24'd247112;
        1767: data_ff <= -24'd131175;
        1768: data_ff <= 24'd71239;
        1769: data_ff <= -24'd37398;
        1770: data_ff <= 24'd18356;
        1771: data_ff <= -24'd8187;
        1772: data_ff <= 24'd3210;
        1773: data_ff <= -24'd1055;
        1774: data_ff <= 24'd266;
        1775: data_ff <= -24'd39;
        1776: data_ff <= 24'd8297247;
        1777: data_ff <= -24'd515079;
        1778: data_ff <= 24'd227370;
        1779: data_ff <= -24'd120279;
        1780: data_ff <= 24'd65116;
        1781: data_ff <= -24'd34078;
        1782: data_ff <= 24'd16673;
        1783: data_ff <= -24'd7412;
        1784: data_ff <= 24'd2896;
        1785: data_ff <= -24'd948;
        1786: data_ff <= 24'd238;
        1787: data_ff <= -24'd35;
        1788: data_ff <= 24'd8309252;
        1789: data_ff <= -24'd472472;
        1790: data_ff <= 24'd207377;
        1791: data_ff <= -24'd109255;
        1792: data_ff <= 24'd58922;
        1793: data_ff <= -24'd30716;
        1794: data_ff <= 24'd14968;
        1795: data_ff <= -24'd6625;
        1796: data_ff <= 24'd2577;
        1797: data_ff <= -24'd840;
        1798: data_ff <= 24'd210;
        1799: data_ff <= -24'd31;
        1800: data_ff <= 24'd8320174;
        1801: data_ff <= -24'd429130;
        1802: data_ff <= 24'd187138;
        1803: data_ff <= -24'd98109;
        1804: data_ff <= 24'd52658;
        1805: data_ff <= -24'd27315;
        1806: data_ff <= 24'd13241;
        1807: data_ff <= -24'd5828;
        1808: data_ff <= 24'd2253;
        1809: data_ff <= -24'd730;
        1810: data_ff <= 24'd181;
        1811: data_ff <= -24'd26;
        1812: data_ff <= 24'd8330012;
        1813: data_ff <= -24'd385057;
        1814: data_ff <= 24'd166660;
        1815: data_ff <= -24'd86842;
        1816: data_ff <= 24'd46328;
        1817: data_ff <= -24'd23876;
        1818: data_ff <= 24'd11493;
        1819: data_ff <= -24'd5020;
        1820: data_ff <= 24'd1925;
        1821: data_ff <= -24'd617;
        1822: data_ff <= 24'd152;
        1823: data_ff <= -24'd22;
        1824: data_ff <= 24'd8338762;
        1825: data_ff <= -24'd340258;
        1826: data_ff <= 24'd145948;
        1827: data_ff <= -24'd75460;
        1828: data_ff <= 24'd39932;
        1829: data_ff <= -24'd20400;
        1830: data_ff <= 24'd9724;
        1831: data_ff <= -24'd4201;
        1832: data_ff <= 24'd1591;
        1833: data_ff <= -24'd503;
        1834: data_ff <= 24'd122;
        1835: data_ff <= -24'd17;
        1836: data_ff <= 24'd8346424;
        1837: data_ff <= -24'd294739;
        1838: data_ff <= 24'd125008;
        1839: data_ff <= -24'd63965;
        1840: data_ff <= 24'd33473;
        1841: data_ff <= -24'd16888;
        1842: data_ff <= 24'd7936;
        1843: data_ff <= -24'd3372;
        1844: data_ff <= 24'd1252;
        1845: data_ff <= -24'd387;
        1846: data_ff <= 24'd91;
        1847: data_ff <= -24'd12;
        1848: data_ff <= 24'd8352994;
        1849: data_ff <= -24'd248506;
        1850: data_ff <= 24'd103847;
        1851: data_ff <= -24'd52361;
        1852: data_ff <= 24'd26953;
        1853: data_ff <= -24'd13341;
        1854: data_ff <= 24'd6129;
        1855: data_ff <= -24'd2534;
        1856: data_ff <= 24'd909;
        1857: data_ff <= -24'd269;
        1858: data_ff <= 24'd60;
        1859: data_ff <= -24'd7;
        1860: data_ff <= 24'd8358472;
        1861: data_ff <= -24'd201564;
        1862: data_ff <= 24'd82471;
        1863: data_ff <= -24'd40652;
        1864: data_ff <= 24'd20374;
        1865: data_ff <= -24'd9760;
        1866: data_ff <= 24'd4302;
        1867: data_ff <= -24'd1685;
        1868: data_ff <= 24'd562;
        1869: data_ff <= -24'd149;
        1870: data_ff <= 24'd28;
        1871: data_ff <= -24'd2;
        1872: data_ff <= 24'd8362856;
        1873: data_ff <= -24'd153919;
        1874: data_ff <= 24'd60886;
        1875: data_ff <= -24'd28842;
        1876: data_ff <= 24'd13739;
        1877: data_ff <= -24'd6147;
        1878: data_ff <= 24'd2458;
        1879: data_ff <= -24'd827;
        1880: data_ff <= 24'd210;
        1881: data_ff <= -24'd27;
        1882: data_ff <= -24'd4;
        1883: data_ff <= 24'd2;
        1884: data_ff <= 24'd8366145;
        1885: data_ff <= -24'd105577;
        1886: data_ff <= 24'd39099;
        1887: data_ff <= -24'd16935;
        1888: data_ff <= 24'd7049;
        1889: data_ff <= -24'd2502;
        1890: data_ff <= 24'd596;
        1891: data_ff <= 24'd39;
        1892: data_ff <= -24'd146;
        1893: data_ff <= 24'd95;
        1894: data_ff <= -24'd37;
        1895: data_ff <= 24'd8;
        1896: data_ff <= 24'd8368338;
        1897: data_ff <= -24'd56546;
        1898: data_ff <= 24'd17116;
        1899: data_ff <= -24'd4935;
        1900: data_ff <= 24'd307;
        1901: data_ff <= 24'd1172;
        1902: data_ff <= -24'd1282;
        1903: data_ff <= 24'd915;
        1904: data_ff <= -24'd507;
        1905: data_ff <= 24'd220;
        1906: data_ff <= -24'd71;
        1907: data_ff <= 24'd13;
        1908: data_ff <= 24'd8369434;
        1909: data_ff <= -24'd6831;
        1910: data_ff <= -24'd5055;
        1911: data_ff <= 24'd7154;
        1912: data_ff <= -24'd6483;
        1913: data_ff <= 24'd4876;
        1914: data_ff <= -24'd3178;
        1915: data_ff <= 24'd1800;
        1916: data_ff <= -24'd872;
        1917: data_ff <= 24'd347;
        1918: data_ff <= -24'd105;
        1919: data_ff <= 24'd19;

        default: data_ff <= 0;
    endcase
end
endmodule
